* Package model for VDD_XLV
* Includes voltage sources and bump connections to M5

* ============================================================================
* Voltage Source for VDD_XLV
* ============================================================================

* Ideal voltage source - value from pg_net_voltage file
v_VDD_XLV VDD_XLV_vsrc 0 VDD_XLV

* ============================================================================
* Bump connections (package rail to M5 die bumps)
* ============================================================================

r VDD_XLV_vsrc VDD_XLV_tap_00000 0.001
r VDD_XLV_tap_00000 8000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00001 0.001
r VDD_XLV_tap_00001 8000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00002 0.001
r VDD_XLV_tap_00002 8000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00003 0.001
r VDD_XLV_tap_00003 8000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00004 0.001
r VDD_XLV_tap_00004 8000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00005 0.001
r VDD_XLV_tap_00005 8000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00006 0.001
r VDD_XLV_tap_00006 8000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00007 0.001
r VDD_XLV_tap_00007 8000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00008 0.001
r VDD_XLV_tap_00008 8000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00009 0.001
r VDD_XLV_tap_00009 8000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00010 0.001
r VDD_XLV_tap_00010 8000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00011 0.001
r VDD_XLV_tap_00011 8000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00012 0.001
r VDD_XLV_tap_00012 16000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00013 0.001
r VDD_XLV_tap_00013 16000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00014 0.001
r VDD_XLV_tap_00014 16000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00015 0.001
r VDD_XLV_tap_00015 16000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00016 0.001
r VDD_XLV_tap_00016 16000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00017 0.001
r VDD_XLV_tap_00017 16000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00018 0.001
r VDD_XLV_tap_00018 16000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00019 0.001
r VDD_XLV_tap_00019 16000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00020 0.001
r VDD_XLV_tap_00020 16000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00021 0.001
r VDD_XLV_tap_00021 16000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00022 0.001
r VDD_XLV_tap_00022 16000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00023 0.001
r VDD_XLV_tap_00023 16000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00024 0.001
r VDD_XLV_tap_00024 24000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00025 0.001
r VDD_XLV_tap_00025 24000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00026 0.001
r VDD_XLV_tap_00026 24000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00027 0.001
r VDD_XLV_tap_00027 24000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00028 0.001
r VDD_XLV_tap_00028 24000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00029 0.001
r VDD_XLV_tap_00029 24000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00030 0.001
r VDD_XLV_tap_00030 24000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00031 0.001
r VDD_XLV_tap_00031 24000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00032 0.001
r VDD_XLV_tap_00032 24000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00033 0.001
r VDD_XLV_tap_00033 24000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00034 0.001
r VDD_XLV_tap_00034 24000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00035 0.001
r VDD_XLV_tap_00035 24000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00036 0.001
r VDD_XLV_tap_00036 32000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00037 0.001
r VDD_XLV_tap_00037 32000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00038 0.001
r VDD_XLV_tap_00038 32000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00039 0.001
r VDD_XLV_tap_00039 32000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00040 0.001
r VDD_XLV_tap_00040 32000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00041 0.001
r VDD_XLV_tap_00041 32000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00042 0.001
r VDD_XLV_tap_00042 32000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00043 0.001
r VDD_XLV_tap_00043 32000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00044 0.001
r VDD_XLV_tap_00044 32000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00045 0.001
r VDD_XLV_tap_00045 32000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00046 0.001
r VDD_XLV_tap_00046 32000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00047 0.001
r VDD_XLV_tap_00047 32000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00048 0.001
r VDD_XLV_tap_00048 40000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00049 0.001
r VDD_XLV_tap_00049 40000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00050 0.001
r VDD_XLV_tap_00050 40000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00051 0.001
r VDD_XLV_tap_00051 40000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00052 0.001
r VDD_XLV_tap_00052 40000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00053 0.001
r VDD_XLV_tap_00053 40000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00054 0.001
r VDD_XLV_tap_00054 40000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00055 0.001
r VDD_XLV_tap_00055 40000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00056 0.001
r VDD_XLV_tap_00056 40000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00057 0.001
r VDD_XLV_tap_00057 40000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00058 0.001
r VDD_XLV_tap_00058 40000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00059 0.001
r VDD_XLV_tap_00059 40000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00060 0.001
r VDD_XLV_tap_00060 48000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00061 0.001
r VDD_XLV_tap_00061 48000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00062 0.001
r VDD_XLV_tap_00062 48000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00063 0.001
r VDD_XLV_tap_00063 48000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00064 0.001
r VDD_XLV_tap_00064 48000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00065 0.001
r VDD_XLV_tap_00065 48000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00066 0.001
r VDD_XLV_tap_00066 48000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00067 0.001
r VDD_XLV_tap_00067 48000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00068 0.001
r VDD_XLV_tap_00068 48000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00069 0.001
r VDD_XLV_tap_00069 48000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00070 0.001
r VDD_XLV_tap_00070 48000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00071 0.001
r VDD_XLV_tap_00071 48000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00072 0.001
r VDD_XLV_tap_00072 56000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00073 0.001
r VDD_XLV_tap_00073 56000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00074 0.001
r VDD_XLV_tap_00074 56000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00075 0.001
r VDD_XLV_tap_00075 56000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00076 0.001
r VDD_XLV_tap_00076 56000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00077 0.001
r VDD_XLV_tap_00077 56000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00078 0.001
r VDD_XLV_tap_00078 56000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00079 0.001
r VDD_XLV_tap_00079 56000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00080 0.001
r VDD_XLV_tap_00080 56000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00081 0.001
r VDD_XLV_tap_00081 56000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00082 0.001
r VDD_XLV_tap_00082 56000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00083 0.001
r VDD_XLV_tap_00083 56000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00084 0.001
r VDD_XLV_tap_00084 64000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00085 0.001
r VDD_XLV_tap_00085 64000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00086 0.001
r VDD_XLV_tap_00086 64000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00087 0.001
r VDD_XLV_tap_00087 64000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00088 0.001
r VDD_XLV_tap_00088 64000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00089 0.001
r VDD_XLV_tap_00089 64000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00090 0.001
r VDD_XLV_tap_00090 64000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00091 0.001
r VDD_XLV_tap_00091 64000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00092 0.001
r VDD_XLV_tap_00092 64000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00093 0.001
r VDD_XLV_tap_00093 64000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00094 0.001
r VDD_XLV_tap_00094 64000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00095 0.001
r VDD_XLV_tap_00095 64000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00096 0.001
r VDD_XLV_tap_00096 72000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00097 0.001
r VDD_XLV_tap_00097 72000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00098 0.001
r VDD_XLV_tap_00098 72000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00099 0.001
r VDD_XLV_tap_00099 72000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00100 0.001
r VDD_XLV_tap_00100 72000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00101 0.001
r VDD_XLV_tap_00101 72000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00102 0.001
r VDD_XLV_tap_00102 72000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00103 0.001
r VDD_XLV_tap_00103 72000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00104 0.001
r VDD_XLV_tap_00104 72000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00105 0.001
r VDD_XLV_tap_00105 72000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00106 0.001
r VDD_XLV_tap_00106 72000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00107 0.001
r VDD_XLV_tap_00107 72000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00108 0.001
r VDD_XLV_tap_00108 80000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00109 0.001
r VDD_XLV_tap_00109 80000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00110 0.001
r VDD_XLV_tap_00110 80000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00111 0.001
r VDD_XLV_tap_00111 80000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00112 0.001
r VDD_XLV_tap_00112 80000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00113 0.001
r VDD_XLV_tap_00113 80000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00114 0.001
r VDD_XLV_tap_00114 80000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00115 0.001
r VDD_XLV_tap_00115 80000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00116 0.001
r VDD_XLV_tap_00116 80000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00117 0.001
r VDD_XLV_tap_00117 80000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00118 0.001
r VDD_XLV_tap_00118 80000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00119 0.001
r VDD_XLV_tap_00119 80000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00120 0.001
r VDD_XLV_tap_00120 88000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00121 0.001
r VDD_XLV_tap_00121 88000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00122 0.001
r VDD_XLV_tap_00122 88000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00123 0.001
r VDD_XLV_tap_00123 88000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00124 0.001
r VDD_XLV_tap_00124 88000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00125 0.001
r VDD_XLV_tap_00125 88000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00126 0.001
r VDD_XLV_tap_00126 88000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00127 0.001
r VDD_XLV_tap_00127 88000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00128 0.001
r VDD_XLV_tap_00128 88000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00129 0.001
r VDD_XLV_tap_00129 88000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00130 0.001
r VDD_XLV_tap_00130 88000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00131 0.001
r VDD_XLV_tap_00131 88000_96000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00132 0.001
r VDD_XLV_tap_00132 96000_8000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00133 0.001
r VDD_XLV_tap_00133 96000_16000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00134 0.001
r VDD_XLV_tap_00134 96000_24000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00135 0.001
r VDD_XLV_tap_00135 96000_32000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00136 0.001
r VDD_XLV_tap_00136 96000_40000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00137 0.001
r VDD_XLV_tap_00137 96000_48000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00138 0.001
r VDD_XLV_tap_00138 96000_56000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00139 0.001
r VDD_XLV_tap_00139 96000_64000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00140 0.001
r VDD_XLV_tap_00140 96000_72000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00141 0.001
r VDD_XLV_tap_00141 96000_80000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00142 0.001
r VDD_XLV_tap_00142 96000_88000_M5 0.001
r VDD_XLV_vsrc VDD_XLV_tap_00143 0.001
r VDD_XLV_tap_00143 96000_96000_M5 0.001