* Tile 0_0 - Die resistor mesh
* 5-layer structure: M1, M2, M3, M4, M5

* ============================================================================
* Layer M1 - 50x50 grid
* ============================================================================

* M1 Horizontal resistors
r 2000_2000_M1 4000_2000_M1 0.020
r 4000_2000_M1 6000_2000_M1 0.020
r 6000_2000_M1 8000_2000_M1 0.020
r 8000_2000_M1 10000_2000_M1 0.020
r 10000_2000_M1 12000_2000_M1 0.020
r 12000_2000_M1 14000_2000_M1 0.020
r 14000_2000_M1 16000_2000_M1 0.020
r 16000_2000_M1 18000_2000_M1 0.020
r 18000_2000_M1 20000_2000_M1 0.020
r 20000_2000_M1 22000_2000_M1 0.020
r 22000_2000_M1 24000_2000_M1 0.020
r 24000_2000_M1 26000_2000_M1 0.020
r 26000_2000_M1 28000_2000_M1 0.020
r 28000_2000_M1 30000_2000_M1 0.020
r 30000_2000_M1 32000_2000_M1 0.020
r 32000_2000_M1 34000_2000_M1 0.020
r 34000_2000_M1 36000_2000_M1 0.020
r 36000_2000_M1 38000_2000_M1 0.020
r 38000_2000_M1 40000_2000_M1 0.020
r 40000_2000_M1 42000_2000_M1 0.020
r 42000_2000_M1 44000_2000_M1 0.020
r 44000_2000_M1 46000_2000_M1 0.020
r 46000_2000_M1 48000_2000_M1 0.020
r 48000_2000_M1 50000_2000_M1 0.020
r 50000_2000_M1 52000_2000_M1 0.020
r 52000_2000_M1 54000_2000_M1 0.020
r 54000_2000_M1 56000_2000_M1 0.020
r 56000_2000_M1 58000_2000_M1 0.020
r 58000_2000_M1 60000_2000_M1 0.020
r 60000_2000_M1 62000_2000_M1 0.020
r 62000_2000_M1 64000_2000_M1 0.020
r 64000_2000_M1 66000_2000_M1 0.020
r 66000_2000_M1 68000_2000_M1 0.020
r 68000_2000_M1 70000_2000_M1 0.020
r 70000_2000_M1 72000_2000_M1 0.020
r 72000_2000_M1 74000_2000_M1 0.020
r 74000_2000_M1 76000_2000_M1 0.020
r 76000_2000_M1 78000_2000_M1 0.020
r 78000_2000_M1 80000_2000_M1 0.020
r 80000_2000_M1 82000_2000_M1 0.020
r 82000_2000_M1 84000_2000_M1 0.020
r 84000_2000_M1 86000_2000_M1 0.020
r 86000_2000_M1 88000_2000_M1 0.020
r 88000_2000_M1 90000_2000_M1 0.020
r 90000_2000_M1 92000_2000_M1 0.020
r 92000_2000_M1 94000_2000_M1 0.020
r 94000_2000_M1 96000_2000_M1 0.020
r 96000_2000_M1 98000_2000_M1 0.020
r 98000_2000_M1 100000_2000_M1 0.020
r 2000_4000_M1 4000_4000_M1 0.020
r 4000_4000_M1 6000_4000_M1 0.020
r 6000_4000_M1 8000_4000_M1 0.020
r 8000_4000_M1 10000_4000_M1 0.020
r 10000_4000_M1 12000_4000_M1 0.020
r 12000_4000_M1 14000_4000_M1 0.020
r 14000_4000_M1 16000_4000_M1 0.020
r 16000_4000_M1 18000_4000_M1 0.020
r 18000_4000_M1 20000_4000_M1 0.020
r 20000_4000_M1 22000_4000_M1 0.020
r 22000_4000_M1 24000_4000_M1 0.020
r 24000_4000_M1 26000_4000_M1 0.020
r 26000_4000_M1 28000_4000_M1 0.020
r 28000_4000_M1 30000_4000_M1 0.020
r 30000_4000_M1 32000_4000_M1 0.020
r 32000_4000_M1 34000_4000_M1 0.020
r 34000_4000_M1 36000_4000_M1 0.020
r 36000_4000_M1 38000_4000_M1 0.020
r 38000_4000_M1 40000_4000_M1 0.020
r 40000_4000_M1 42000_4000_M1 0.020
r 42000_4000_M1 44000_4000_M1 0.020
r 44000_4000_M1 46000_4000_M1 0.020
r 46000_4000_M1 48000_4000_M1 0.020
r 48000_4000_M1 50000_4000_M1 0.020
r 50000_4000_M1 52000_4000_M1 0.020
r 52000_4000_M1 54000_4000_M1 0.020
r 54000_4000_M1 56000_4000_M1 0.020
r 56000_4000_M1 58000_4000_M1 0.020
r 58000_4000_M1 60000_4000_M1 0.020
r 60000_4000_M1 62000_4000_M1 0.020
r 62000_4000_M1 64000_4000_M1 0.020
r 64000_4000_M1 66000_4000_M1 0.020
r 66000_4000_M1 68000_4000_M1 0.020
r 68000_4000_M1 70000_4000_M1 0.020
r 70000_4000_M1 72000_4000_M1 0.020
r 72000_4000_M1 74000_4000_M1 0.020
r 74000_4000_M1 76000_4000_M1 0.020
r 76000_4000_M1 78000_4000_M1 0.020
r 78000_4000_M1 80000_4000_M1 0.020
r 80000_4000_M1 82000_4000_M1 0.020
r 82000_4000_M1 84000_4000_M1 0.020
r 84000_4000_M1 86000_4000_M1 0.020
r 86000_4000_M1 88000_4000_M1 0.020
r 88000_4000_M1 90000_4000_M1 0.020
r 90000_4000_M1 92000_4000_M1 0.020
r 92000_4000_M1 94000_4000_M1 0.020
r 94000_4000_M1 96000_4000_M1 0.020
r 96000_4000_M1 98000_4000_M1 0.020
r 98000_4000_M1 100000_4000_M1 0.020
r 2000_6000_M1 4000_6000_M1 0.020
r 4000_6000_M1 6000_6000_M1 0.020
r 6000_6000_M1 8000_6000_M1 0.020
r 8000_6000_M1 10000_6000_M1 0.020
r 10000_6000_M1 12000_6000_M1 0.020
r 12000_6000_M1 14000_6000_M1 0.020
r 14000_6000_M1 16000_6000_M1 0.020
r 16000_6000_M1 18000_6000_M1 0.020
r 18000_6000_M1 20000_6000_M1 0.020
r 20000_6000_M1 22000_6000_M1 0.020
r 22000_6000_M1 24000_6000_M1 0.020
r 24000_6000_M1 26000_6000_M1 0.020
r 26000_6000_M1 28000_6000_M1 0.020
r 28000_6000_M1 30000_6000_M1 0.020
r 30000_6000_M1 32000_6000_M1 0.020
r 32000_6000_M1 34000_6000_M1 0.020
r 34000_6000_M1 36000_6000_M1 0.020
r 36000_6000_M1 38000_6000_M1 0.020
r 38000_6000_M1 40000_6000_M1 0.020
r 40000_6000_M1 42000_6000_M1 0.020
r 42000_6000_M1 44000_6000_M1 0.020
r 44000_6000_M1 46000_6000_M1 0.020
r 46000_6000_M1 48000_6000_M1 0.020
r 48000_6000_M1 50000_6000_M1 0.020
r 50000_6000_M1 52000_6000_M1 0.020
r 52000_6000_M1 54000_6000_M1 0.020
r 54000_6000_M1 56000_6000_M1 0.020
r 56000_6000_M1 58000_6000_M1 0.020
r 58000_6000_M1 60000_6000_M1 0.020
r 60000_6000_M1 62000_6000_M1 0.020
r 62000_6000_M1 64000_6000_M1 0.020
r 64000_6000_M1 66000_6000_M1 0.020
r 66000_6000_M1 68000_6000_M1 0.020
r 68000_6000_M1 70000_6000_M1 0.020
r 70000_6000_M1 72000_6000_M1 0.020
r 72000_6000_M1 74000_6000_M1 0.020
r 74000_6000_M1 76000_6000_M1 0.020
r 76000_6000_M1 78000_6000_M1 0.020
r 78000_6000_M1 80000_6000_M1 0.020
r 80000_6000_M1 82000_6000_M1 0.020
r 82000_6000_M1 84000_6000_M1 0.020
r 84000_6000_M1 86000_6000_M1 0.020
r 86000_6000_M1 88000_6000_M1 0.020
r 88000_6000_M1 90000_6000_M1 0.020
r 90000_6000_M1 92000_6000_M1 0.020
r 92000_6000_M1 94000_6000_M1 0.020
r 94000_6000_M1 96000_6000_M1 0.020
r 96000_6000_M1 98000_6000_M1 0.020
r 98000_6000_M1 100000_6000_M1 0.020
r 2000_8000_M1 4000_8000_M1 0.020
r 4000_8000_M1 6000_8000_M1 0.020
r 6000_8000_M1 8000_8000_M1 0.020
r 8000_8000_M1 10000_8000_M1 0.020
r 10000_8000_M1 12000_8000_M1 0.020
r 12000_8000_M1 14000_8000_M1 0.020
r 14000_8000_M1 16000_8000_M1 0.020
r 16000_8000_M1 18000_8000_M1 0.020
r 18000_8000_M1 20000_8000_M1 0.020
r 20000_8000_M1 22000_8000_M1 0.020
r 22000_8000_M1 24000_8000_M1 0.020
r 24000_8000_M1 26000_8000_M1 0.020
r 26000_8000_M1 28000_8000_M1 0.020
r 28000_8000_M1 30000_8000_M1 0.020
r 30000_8000_M1 32000_8000_M1 0.020
r 32000_8000_M1 34000_8000_M1 0.020
r 34000_8000_M1 36000_8000_M1 0.020
r 36000_8000_M1 38000_8000_M1 0.020
r 38000_8000_M1 40000_8000_M1 0.020
r 40000_8000_M1 42000_8000_M1 0.020
r 42000_8000_M1 44000_8000_M1 0.020
r 44000_8000_M1 46000_8000_M1 0.020
r 46000_8000_M1 48000_8000_M1 0.020
r 48000_8000_M1 50000_8000_M1 0.020
r 50000_8000_M1 52000_8000_M1 0.020
r 52000_8000_M1 54000_8000_M1 0.020
r 54000_8000_M1 56000_8000_M1 0.020
r 56000_8000_M1 58000_8000_M1 0.020
r 58000_8000_M1 60000_8000_M1 0.020
r 60000_8000_M1 62000_8000_M1 0.020
r 62000_8000_M1 64000_8000_M1 0.020
r 64000_8000_M1 66000_8000_M1 0.020
r 66000_8000_M1 68000_8000_M1 0.020
r 68000_8000_M1 70000_8000_M1 0.020
r 70000_8000_M1 72000_8000_M1 0.020
r 72000_8000_M1 74000_8000_M1 0.020
r 74000_8000_M1 76000_8000_M1 0.020
r 76000_8000_M1 78000_8000_M1 0.020
r 78000_8000_M1 80000_8000_M1 0.020
r 80000_8000_M1 82000_8000_M1 0.020
r 82000_8000_M1 84000_8000_M1 0.020
r 84000_8000_M1 86000_8000_M1 0.020
r 86000_8000_M1 88000_8000_M1 0.020
r 88000_8000_M1 90000_8000_M1 0.020
r 90000_8000_M1 92000_8000_M1 0.020
r 92000_8000_M1 94000_8000_M1 0.020
r 94000_8000_M1 96000_8000_M1 0.020
r 96000_8000_M1 98000_8000_M1 0.020
r 98000_8000_M1 100000_8000_M1 0.020
r 2000_10000_M1 4000_10000_M1 0.020
r 4000_10000_M1 6000_10000_M1 0.020
r 6000_10000_M1 8000_10000_M1 0.020
r 8000_10000_M1 10000_10000_M1 0.020
r 10000_10000_M1 12000_10000_M1 0.020
r 12000_10000_M1 14000_10000_M1 0.020
r 14000_10000_M1 16000_10000_M1 0.020
r 16000_10000_M1 18000_10000_M1 0.020
r 18000_10000_M1 20000_10000_M1 0.020
r 20000_10000_M1 22000_10000_M1 0.020
r 22000_10000_M1 24000_10000_M1 0.020
r 24000_10000_M1 26000_10000_M1 0.020
r 26000_10000_M1 28000_10000_M1 0.020
r 28000_10000_M1 30000_10000_M1 0.020
r 30000_10000_M1 32000_10000_M1 0.020
r 32000_10000_M1 34000_10000_M1 0.020
r 34000_10000_M1 36000_10000_M1 0.020
r 36000_10000_M1 38000_10000_M1 0.020
r 38000_10000_M1 40000_10000_M1 0.020
r 40000_10000_M1 42000_10000_M1 0.020
r 42000_10000_M1 44000_10000_M1 0.020
r 44000_10000_M1 46000_10000_M1 0.020
r 46000_10000_M1 48000_10000_M1 0.020
r 48000_10000_M1 50000_10000_M1 0.020
r 50000_10000_M1 52000_10000_M1 0.020
r 52000_10000_M1 54000_10000_M1 0.020
r 54000_10000_M1 56000_10000_M1 0.020
r 56000_10000_M1 58000_10000_M1 0.020
r 58000_10000_M1 60000_10000_M1 0.020
r 60000_10000_M1 62000_10000_M1 0.020
r 62000_10000_M1 64000_10000_M1 0.020
r 64000_10000_M1 66000_10000_M1 0.020
r 66000_10000_M1 68000_10000_M1 0.020
r 68000_10000_M1 70000_10000_M1 0.020
r 70000_10000_M1 72000_10000_M1 0.020
r 72000_10000_M1 74000_10000_M1 0.020
r 74000_10000_M1 76000_10000_M1 0.020
r 76000_10000_M1 78000_10000_M1 0.020
r 78000_10000_M1 80000_10000_M1 0.020
r 80000_10000_M1 82000_10000_M1 0.020
r 82000_10000_M1 84000_10000_M1 0.020
r 84000_10000_M1 86000_10000_M1 0.020
r 86000_10000_M1 88000_10000_M1 0.020
r 88000_10000_M1 90000_10000_M1 0.020
r 90000_10000_M1 92000_10000_M1 0.020
r 92000_10000_M1 94000_10000_M1 0.020
r 94000_10000_M1 96000_10000_M1 0.020
r 96000_10000_M1 98000_10000_M1 0.020
r 98000_10000_M1 100000_10000_M1 0.020
r 2000_12000_M1 4000_12000_M1 0.020
r 4000_12000_M1 6000_12000_M1 0.020
r 6000_12000_M1 8000_12000_M1 0.020
r 8000_12000_M1 10000_12000_M1 0.020
r 10000_12000_M1 12000_12000_M1 0.020
r 12000_12000_M1 14000_12000_M1 0.020
r 14000_12000_M1 16000_12000_M1 0.020
r 16000_12000_M1 18000_12000_M1 0.020
r 18000_12000_M1 20000_12000_M1 0.020
r 20000_12000_M1 22000_12000_M1 0.020
r 22000_12000_M1 24000_12000_M1 0.020
r 24000_12000_M1 26000_12000_M1 0.020
r 26000_12000_M1 28000_12000_M1 0.020
r 28000_12000_M1 30000_12000_M1 0.020
r 30000_12000_M1 32000_12000_M1 0.020
r 32000_12000_M1 34000_12000_M1 0.020
r 34000_12000_M1 36000_12000_M1 0.020
r 36000_12000_M1 38000_12000_M1 0.020
r 38000_12000_M1 40000_12000_M1 0.020
r 40000_12000_M1 42000_12000_M1 0.020
r 42000_12000_M1 44000_12000_M1 0.020
r 44000_12000_M1 46000_12000_M1 0.020
r 46000_12000_M1 48000_12000_M1 0.020
r 48000_12000_M1 50000_12000_M1 0.020
r 50000_12000_M1 52000_12000_M1 0.020
r 52000_12000_M1 54000_12000_M1 0.020
r 54000_12000_M1 56000_12000_M1 0.020
r 56000_12000_M1 58000_12000_M1 0.020
r 58000_12000_M1 60000_12000_M1 0.020
r 60000_12000_M1 62000_12000_M1 0.020
r 62000_12000_M1 64000_12000_M1 0.020
r 64000_12000_M1 66000_12000_M1 0.020
r 66000_12000_M1 68000_12000_M1 0.020
r 68000_12000_M1 70000_12000_M1 0.020
r 70000_12000_M1 72000_12000_M1 0.020
r 72000_12000_M1 74000_12000_M1 0.020
r 74000_12000_M1 76000_12000_M1 0.020
r 76000_12000_M1 78000_12000_M1 0.020
r 78000_12000_M1 80000_12000_M1 0.020
r 80000_12000_M1 82000_12000_M1 0.020
r 82000_12000_M1 84000_12000_M1 0.020
r 84000_12000_M1 86000_12000_M1 0.020
r 86000_12000_M1 88000_12000_M1 0.020
r 88000_12000_M1 90000_12000_M1 0.020
r 90000_12000_M1 92000_12000_M1 0.020
r 92000_12000_M1 94000_12000_M1 0.020
r 94000_12000_M1 96000_12000_M1 0.020
r 96000_12000_M1 98000_12000_M1 0.020
r 98000_12000_M1 100000_12000_M1 0.020
r 2000_14000_M1 4000_14000_M1 0.020
r 4000_14000_M1 6000_14000_M1 0.020
r 6000_14000_M1 8000_14000_M1 0.020
r 8000_14000_M1 10000_14000_M1 0.020
r 10000_14000_M1 12000_14000_M1 0.020
r 12000_14000_M1 14000_14000_M1 0.020
r 14000_14000_M1 16000_14000_M1 0.020
r 16000_14000_M1 18000_14000_M1 0.020
r 18000_14000_M1 20000_14000_M1 0.020
r 20000_14000_M1 22000_14000_M1 0.020
r 22000_14000_M1 24000_14000_M1 0.020
r 24000_14000_M1 26000_14000_M1 0.020
r 26000_14000_M1 28000_14000_M1 0.020
r 28000_14000_M1 30000_14000_M1 0.020
r 30000_14000_M1 32000_14000_M1 0.020
r 32000_14000_M1 34000_14000_M1 0.020
r 34000_14000_M1 36000_14000_M1 0.020
r 36000_14000_M1 38000_14000_M1 0.020
r 38000_14000_M1 40000_14000_M1 0.020
r 40000_14000_M1 42000_14000_M1 0.020
r 42000_14000_M1 44000_14000_M1 0.020
r 44000_14000_M1 46000_14000_M1 0.020
r 46000_14000_M1 48000_14000_M1 0.020
r 48000_14000_M1 50000_14000_M1 0.020
r 50000_14000_M1 52000_14000_M1 0.020
r 52000_14000_M1 54000_14000_M1 0.020
r 54000_14000_M1 56000_14000_M1 0.020
r 56000_14000_M1 58000_14000_M1 0.020
r 58000_14000_M1 60000_14000_M1 0.020
r 60000_14000_M1 62000_14000_M1 0.020
r 62000_14000_M1 64000_14000_M1 0.020
r 64000_14000_M1 66000_14000_M1 0.020
r 66000_14000_M1 68000_14000_M1 0.020
r 68000_14000_M1 70000_14000_M1 0.020
r 70000_14000_M1 72000_14000_M1 0.020
r 72000_14000_M1 74000_14000_M1 0.020
r 74000_14000_M1 76000_14000_M1 0.020
r 76000_14000_M1 78000_14000_M1 0.020
r 78000_14000_M1 80000_14000_M1 0.020
r 80000_14000_M1 82000_14000_M1 0.020
r 82000_14000_M1 84000_14000_M1 0.020
r 84000_14000_M1 86000_14000_M1 0.020
r 86000_14000_M1 88000_14000_M1 0.020
r 88000_14000_M1 90000_14000_M1 0.020
r 90000_14000_M1 92000_14000_M1 0.020
r 92000_14000_M1 94000_14000_M1 0.020
r 94000_14000_M1 96000_14000_M1 0.020
r 96000_14000_M1 98000_14000_M1 0.020
r 98000_14000_M1 100000_14000_M1 0.020
r 2000_16000_M1 4000_16000_M1 0.020
r 4000_16000_M1 6000_16000_M1 0.020
r 6000_16000_M1 8000_16000_M1 0.020
r 8000_16000_M1 10000_16000_M1 0.020
r 10000_16000_M1 12000_16000_M1 0.020
r 12000_16000_M1 14000_16000_M1 0.020
r 14000_16000_M1 16000_16000_M1 0.020
r 16000_16000_M1 18000_16000_M1 0.020
r 18000_16000_M1 20000_16000_M1 0.020
r 20000_16000_M1 22000_16000_M1 0.020
r 22000_16000_M1 24000_16000_M1 0.020
r 24000_16000_M1 26000_16000_M1 0.020
r 26000_16000_M1 28000_16000_M1 0.020
r 28000_16000_M1 30000_16000_M1 0.020
r 30000_16000_M1 32000_16000_M1 0.020
r 32000_16000_M1 34000_16000_M1 0.020
r 34000_16000_M1 36000_16000_M1 0.020
r 36000_16000_M1 38000_16000_M1 0.020
r 38000_16000_M1 40000_16000_M1 0.020
r 40000_16000_M1 42000_16000_M1 0.020
r 42000_16000_M1 44000_16000_M1 0.020
r 44000_16000_M1 46000_16000_M1 0.020
r 46000_16000_M1 48000_16000_M1 0.020
r 48000_16000_M1 50000_16000_M1 0.020
r 50000_16000_M1 52000_16000_M1 0.020
r 52000_16000_M1 54000_16000_M1 0.020
r 54000_16000_M1 56000_16000_M1 0.020
r 56000_16000_M1 58000_16000_M1 0.020
r 58000_16000_M1 60000_16000_M1 0.020
r 60000_16000_M1 62000_16000_M1 0.020
r 62000_16000_M1 64000_16000_M1 0.020
r 64000_16000_M1 66000_16000_M1 0.020
r 66000_16000_M1 68000_16000_M1 0.020
r 68000_16000_M1 70000_16000_M1 0.020
r 70000_16000_M1 72000_16000_M1 0.020
r 72000_16000_M1 74000_16000_M1 0.020
r 74000_16000_M1 76000_16000_M1 0.020
r 76000_16000_M1 78000_16000_M1 0.020
r 78000_16000_M1 80000_16000_M1 0.020
r 80000_16000_M1 82000_16000_M1 0.020
r 82000_16000_M1 84000_16000_M1 0.020
r 84000_16000_M1 86000_16000_M1 0.020
r 86000_16000_M1 88000_16000_M1 0.020
r 88000_16000_M1 90000_16000_M1 0.020
r 90000_16000_M1 92000_16000_M1 0.020
r 92000_16000_M1 94000_16000_M1 0.020
r 94000_16000_M1 96000_16000_M1 0.020
r 96000_16000_M1 98000_16000_M1 0.020
r 98000_16000_M1 100000_16000_M1 0.020
r 2000_18000_M1 4000_18000_M1 0.020
r 4000_18000_M1 6000_18000_M1 0.020
r 6000_18000_M1 8000_18000_M1 0.020
r 8000_18000_M1 10000_18000_M1 0.020
r 10000_18000_M1 12000_18000_M1 0.020
r 12000_18000_M1 14000_18000_M1 0.020
r 14000_18000_M1 16000_18000_M1 0.020
r 16000_18000_M1 18000_18000_M1 0.020
r 18000_18000_M1 20000_18000_M1 0.020
r 20000_18000_M1 22000_18000_M1 0.020
r 22000_18000_M1 24000_18000_M1 0.020
r 24000_18000_M1 26000_18000_M1 0.020
r 26000_18000_M1 28000_18000_M1 0.020
r 28000_18000_M1 30000_18000_M1 0.020
r 30000_18000_M1 32000_18000_M1 0.020
r 32000_18000_M1 34000_18000_M1 0.020
r 34000_18000_M1 36000_18000_M1 0.020
r 36000_18000_M1 38000_18000_M1 0.020
r 38000_18000_M1 40000_18000_M1 0.020
r 40000_18000_M1 42000_18000_M1 0.020
r 42000_18000_M1 44000_18000_M1 0.020
r 44000_18000_M1 46000_18000_M1 0.020
r 46000_18000_M1 48000_18000_M1 0.020
r 48000_18000_M1 50000_18000_M1 0.020
r 50000_18000_M1 52000_18000_M1 0.020
r 52000_18000_M1 54000_18000_M1 0.020
r 54000_18000_M1 56000_18000_M1 0.020
r 56000_18000_M1 58000_18000_M1 0.020
r 58000_18000_M1 60000_18000_M1 0.020
r 60000_18000_M1 62000_18000_M1 0.020
r 62000_18000_M1 64000_18000_M1 0.020
r 64000_18000_M1 66000_18000_M1 0.020
r 66000_18000_M1 68000_18000_M1 0.020
r 68000_18000_M1 70000_18000_M1 0.020
r 70000_18000_M1 72000_18000_M1 0.020
r 72000_18000_M1 74000_18000_M1 0.020
r 74000_18000_M1 76000_18000_M1 0.020
r 76000_18000_M1 78000_18000_M1 0.020
r 78000_18000_M1 80000_18000_M1 0.020
r 80000_18000_M1 82000_18000_M1 0.020
r 82000_18000_M1 84000_18000_M1 0.020
r 84000_18000_M1 86000_18000_M1 0.020
r 86000_18000_M1 88000_18000_M1 0.020
r 88000_18000_M1 90000_18000_M1 0.020
r 90000_18000_M1 92000_18000_M1 0.020
r 92000_18000_M1 94000_18000_M1 0.020
r 94000_18000_M1 96000_18000_M1 0.020
r 96000_18000_M1 98000_18000_M1 0.020
r 98000_18000_M1 100000_18000_M1 0.020
r 2000_20000_M1 4000_20000_M1 0.020
r 4000_20000_M1 6000_20000_M1 0.020
r 6000_20000_M1 8000_20000_M1 0.020
r 8000_20000_M1 10000_20000_M1 0.020
r 10000_20000_M1 12000_20000_M1 0.020
r 12000_20000_M1 14000_20000_M1 0.020
r 14000_20000_M1 16000_20000_M1 0.020
r 16000_20000_M1 18000_20000_M1 0.020
r 18000_20000_M1 20000_20000_M1 0.020
r 20000_20000_M1 22000_20000_M1 0.020
r 22000_20000_M1 24000_20000_M1 0.020
r 24000_20000_M1 26000_20000_M1 0.020
r 26000_20000_M1 28000_20000_M1 0.020
r 28000_20000_M1 30000_20000_M1 0.020
r 30000_20000_M1 32000_20000_M1 0.020
r 32000_20000_M1 34000_20000_M1 0.020
r 34000_20000_M1 36000_20000_M1 0.020
r 36000_20000_M1 38000_20000_M1 0.020
r 38000_20000_M1 40000_20000_M1 0.020
r 40000_20000_M1 42000_20000_M1 0.020
r 42000_20000_M1 44000_20000_M1 0.020
r 44000_20000_M1 46000_20000_M1 0.020
r 46000_20000_M1 48000_20000_M1 0.020
r 48000_20000_M1 50000_20000_M1 0.020
r 50000_20000_M1 52000_20000_M1 0.020
r 52000_20000_M1 54000_20000_M1 0.020
r 54000_20000_M1 56000_20000_M1 0.020
r 56000_20000_M1 58000_20000_M1 0.020
r 58000_20000_M1 60000_20000_M1 0.020
r 60000_20000_M1 62000_20000_M1 0.020
r 62000_20000_M1 64000_20000_M1 0.020
r 64000_20000_M1 66000_20000_M1 0.020
r 66000_20000_M1 68000_20000_M1 0.020
r 68000_20000_M1 70000_20000_M1 0.020
r 70000_20000_M1 72000_20000_M1 0.020
r 72000_20000_M1 74000_20000_M1 0.020
r 74000_20000_M1 76000_20000_M1 0.020
r 76000_20000_M1 78000_20000_M1 0.020
r 78000_20000_M1 80000_20000_M1 0.020
r 80000_20000_M1 82000_20000_M1 0.020
r 82000_20000_M1 84000_20000_M1 0.020
r 84000_20000_M1 86000_20000_M1 0.020
r 86000_20000_M1 88000_20000_M1 0.020
r 88000_20000_M1 90000_20000_M1 0.020
r 90000_20000_M1 92000_20000_M1 0.020
r 92000_20000_M1 94000_20000_M1 0.020
r 94000_20000_M1 96000_20000_M1 0.020
r 96000_20000_M1 98000_20000_M1 0.020
r 98000_20000_M1 100000_20000_M1 0.020
r 2000_22000_M1 4000_22000_M1 0.020
r 4000_22000_M1 6000_22000_M1 0.020
r 6000_22000_M1 8000_22000_M1 0.020
r 8000_22000_M1 10000_22000_M1 0.020
r 10000_22000_M1 12000_22000_M1 0.020
r 12000_22000_M1 14000_22000_M1 0.020
r 14000_22000_M1 16000_22000_M1 0.020
r 16000_22000_M1 18000_22000_M1 0.020
r 18000_22000_M1 20000_22000_M1 0.020
r 20000_22000_M1 22000_22000_M1 0.020
r 22000_22000_M1 24000_22000_M1 0.020
r 24000_22000_M1 26000_22000_M1 0.020
r 26000_22000_M1 28000_22000_M1 0.020
r 28000_22000_M1 30000_22000_M1 0.020
r 30000_22000_M1 32000_22000_M1 0.020
r 32000_22000_M1 34000_22000_M1 0.020
r 34000_22000_M1 36000_22000_M1 0.020
r 36000_22000_M1 38000_22000_M1 0.020
r 38000_22000_M1 40000_22000_M1 0.020
r 40000_22000_M1 42000_22000_M1 0.020
r 42000_22000_M1 44000_22000_M1 0.020
r 44000_22000_M1 46000_22000_M1 0.020
r 46000_22000_M1 48000_22000_M1 0.020
r 48000_22000_M1 50000_22000_M1 0.020
r 50000_22000_M1 52000_22000_M1 0.020
r 52000_22000_M1 54000_22000_M1 0.020
r 54000_22000_M1 56000_22000_M1 0.020
r 56000_22000_M1 58000_22000_M1 0.020
r 58000_22000_M1 60000_22000_M1 0.020
r 60000_22000_M1 62000_22000_M1 0.020
r 62000_22000_M1 64000_22000_M1 0.020
r 64000_22000_M1 66000_22000_M1 0.020
r 66000_22000_M1 68000_22000_M1 0.020
r 68000_22000_M1 70000_22000_M1 0.020
r 70000_22000_M1 72000_22000_M1 0.020
r 72000_22000_M1 74000_22000_M1 0.020
r 74000_22000_M1 76000_22000_M1 0.020
r 76000_22000_M1 78000_22000_M1 0.020
r 78000_22000_M1 80000_22000_M1 0.020
r 80000_22000_M1 82000_22000_M1 0.020
r 82000_22000_M1 84000_22000_M1 0.020
r 84000_22000_M1 86000_22000_M1 0.020
r 86000_22000_M1 88000_22000_M1 0.020
r 88000_22000_M1 90000_22000_M1 0.020
r 90000_22000_M1 92000_22000_M1 0.020
r 92000_22000_M1 94000_22000_M1 0.020
r 94000_22000_M1 96000_22000_M1 0.020
r 96000_22000_M1 98000_22000_M1 0.020
r 98000_22000_M1 100000_22000_M1 0.020
r 2000_24000_M1 4000_24000_M1 0.020
r 4000_24000_M1 6000_24000_M1 0.020
r 6000_24000_M1 8000_24000_M1 0.020
r 8000_24000_M1 10000_24000_M1 0.020
r 10000_24000_M1 12000_24000_M1 0.020
r 12000_24000_M1 14000_24000_M1 0.020
r 14000_24000_M1 16000_24000_M1 0.020
r 16000_24000_M1 18000_24000_M1 0.020
r 18000_24000_M1 20000_24000_M1 0.020
r 20000_24000_M1 22000_24000_M1 0.020
r 22000_24000_M1 24000_24000_M1 0.020
r 24000_24000_M1 26000_24000_M1 0.020
r 26000_24000_M1 28000_24000_M1 0.020
r 28000_24000_M1 30000_24000_M1 0.020
r 30000_24000_M1 32000_24000_M1 0.020
r 32000_24000_M1 34000_24000_M1 0.020
r 34000_24000_M1 36000_24000_M1 0.020
r 36000_24000_M1 38000_24000_M1 0.020
r 38000_24000_M1 40000_24000_M1 0.020
r 40000_24000_M1 42000_24000_M1 0.020
r 42000_24000_M1 44000_24000_M1 0.020
r 44000_24000_M1 46000_24000_M1 0.020
r 46000_24000_M1 48000_24000_M1 0.020
r 48000_24000_M1 50000_24000_M1 0.020
r 50000_24000_M1 52000_24000_M1 0.020
r 52000_24000_M1 54000_24000_M1 0.020
r 54000_24000_M1 56000_24000_M1 0.020
r 56000_24000_M1 58000_24000_M1 0.020
r 58000_24000_M1 60000_24000_M1 0.020
r 60000_24000_M1 62000_24000_M1 0.020
r 62000_24000_M1 64000_24000_M1 0.020
r 64000_24000_M1 66000_24000_M1 0.020
r 66000_24000_M1 68000_24000_M1 0.020
r 68000_24000_M1 70000_24000_M1 0.020
r 70000_24000_M1 72000_24000_M1 0.020
r 72000_24000_M1 74000_24000_M1 0.020
r 74000_24000_M1 76000_24000_M1 0.020
r 76000_24000_M1 78000_24000_M1 0.020
r 78000_24000_M1 80000_24000_M1 0.020
r 80000_24000_M1 82000_24000_M1 0.020
r 82000_24000_M1 84000_24000_M1 0.020
r 84000_24000_M1 86000_24000_M1 0.020
r 86000_24000_M1 88000_24000_M1 0.020
r 88000_24000_M1 90000_24000_M1 0.020
r 90000_24000_M1 92000_24000_M1 0.020
r 92000_24000_M1 94000_24000_M1 0.020
r 94000_24000_M1 96000_24000_M1 0.020
r 96000_24000_M1 98000_24000_M1 0.020
r 98000_24000_M1 100000_24000_M1 0.020
r 2000_26000_M1 4000_26000_M1 0.020
r 4000_26000_M1 6000_26000_M1 0.020
r 6000_26000_M1 8000_26000_M1 0.020
r 8000_26000_M1 10000_26000_M1 0.020
r 10000_26000_M1 12000_26000_M1 0.020
r 12000_26000_M1 14000_26000_M1 0.020
r 14000_26000_M1 16000_26000_M1 0.020
r 16000_26000_M1 18000_26000_M1 0.020
r 18000_26000_M1 20000_26000_M1 0.020
r 20000_26000_M1 22000_26000_M1 0.020
r 22000_26000_M1 24000_26000_M1 0.020
r 24000_26000_M1 26000_26000_M1 0.020
r 26000_26000_M1 28000_26000_M1 0.020
r 28000_26000_M1 30000_26000_M1 0.020
r 30000_26000_M1 32000_26000_M1 0.020
r 32000_26000_M1 34000_26000_M1 0.020
r 34000_26000_M1 36000_26000_M1 0.020
r 36000_26000_M1 38000_26000_M1 0.020
r 38000_26000_M1 40000_26000_M1 0.020
r 40000_26000_M1 42000_26000_M1 0.020
r 42000_26000_M1 44000_26000_M1 0.020
r 44000_26000_M1 46000_26000_M1 0.020
r 46000_26000_M1 48000_26000_M1 0.020
r 48000_26000_M1 50000_26000_M1 0.020
r 50000_26000_M1 52000_26000_M1 0.020
r 52000_26000_M1 54000_26000_M1 0.020
r 54000_26000_M1 56000_26000_M1 0.020
r 56000_26000_M1 58000_26000_M1 0.020
r 58000_26000_M1 60000_26000_M1 0.020
r 60000_26000_M1 62000_26000_M1 0.020
r 62000_26000_M1 64000_26000_M1 0.020
r 64000_26000_M1 66000_26000_M1 0.020
r 66000_26000_M1 68000_26000_M1 0.020
r 68000_26000_M1 70000_26000_M1 0.020
r 70000_26000_M1 72000_26000_M1 0.020
r 72000_26000_M1 74000_26000_M1 0.020
r 74000_26000_M1 76000_26000_M1 0.020
r 76000_26000_M1 78000_26000_M1 0.020
r 78000_26000_M1 80000_26000_M1 0.020
r 80000_26000_M1 82000_26000_M1 0.020
r 82000_26000_M1 84000_26000_M1 0.020
r 84000_26000_M1 86000_26000_M1 0.020
r 86000_26000_M1 88000_26000_M1 0.020
r 88000_26000_M1 90000_26000_M1 0.020
r 90000_26000_M1 92000_26000_M1 0.020
r 92000_26000_M1 94000_26000_M1 0.020
r 94000_26000_M1 96000_26000_M1 0.020
r 96000_26000_M1 98000_26000_M1 0.020
r 98000_26000_M1 100000_26000_M1 0.020
r 2000_28000_M1 4000_28000_M1 0.020
r 4000_28000_M1 6000_28000_M1 0.020
r 6000_28000_M1 8000_28000_M1 0.020
r 8000_28000_M1 10000_28000_M1 0.020
r 10000_28000_M1 12000_28000_M1 0.020
r 12000_28000_M1 14000_28000_M1 0.020
r 14000_28000_M1 16000_28000_M1 0.020
r 16000_28000_M1 18000_28000_M1 0.020
r 18000_28000_M1 20000_28000_M1 0.020
r 20000_28000_M1 22000_28000_M1 0.020
r 22000_28000_M1 24000_28000_M1 0.020
r 24000_28000_M1 26000_28000_M1 0.020
r 26000_28000_M1 28000_28000_M1 0.020
r 28000_28000_M1 30000_28000_M1 0.020
r 30000_28000_M1 32000_28000_M1 0.020
r 32000_28000_M1 34000_28000_M1 0.020
r 34000_28000_M1 36000_28000_M1 0.020
r 36000_28000_M1 38000_28000_M1 0.020
r 38000_28000_M1 40000_28000_M1 0.020
r 40000_28000_M1 42000_28000_M1 0.020
r 42000_28000_M1 44000_28000_M1 0.020
r 44000_28000_M1 46000_28000_M1 0.020
r 46000_28000_M1 48000_28000_M1 0.020
r 48000_28000_M1 50000_28000_M1 0.020
r 50000_28000_M1 52000_28000_M1 0.020
r 52000_28000_M1 54000_28000_M1 0.020
r 54000_28000_M1 56000_28000_M1 0.020
r 56000_28000_M1 58000_28000_M1 0.020
r 58000_28000_M1 60000_28000_M1 0.020
r 60000_28000_M1 62000_28000_M1 0.020
r 62000_28000_M1 64000_28000_M1 0.020
r 64000_28000_M1 66000_28000_M1 0.020
r 66000_28000_M1 68000_28000_M1 0.020
r 68000_28000_M1 70000_28000_M1 0.020
r 70000_28000_M1 72000_28000_M1 0.020
r 72000_28000_M1 74000_28000_M1 0.020
r 74000_28000_M1 76000_28000_M1 0.020
r 76000_28000_M1 78000_28000_M1 0.020
r 78000_28000_M1 80000_28000_M1 0.020
r 80000_28000_M1 82000_28000_M1 0.020
r 82000_28000_M1 84000_28000_M1 0.020
r 84000_28000_M1 86000_28000_M1 0.020
r 86000_28000_M1 88000_28000_M1 0.020
r 88000_28000_M1 90000_28000_M1 0.020
r 90000_28000_M1 92000_28000_M1 0.020
r 92000_28000_M1 94000_28000_M1 0.020
r 94000_28000_M1 96000_28000_M1 0.020
r 96000_28000_M1 98000_28000_M1 0.020
r 98000_28000_M1 100000_28000_M1 0.020
r 2000_30000_M1 4000_30000_M1 0.020
r 4000_30000_M1 6000_30000_M1 0.020
r 6000_30000_M1 8000_30000_M1 0.020
r 8000_30000_M1 10000_30000_M1 0.020
r 10000_30000_M1 12000_30000_M1 0.020
r 12000_30000_M1 14000_30000_M1 0.020
r 14000_30000_M1 16000_30000_M1 0.020
r 16000_30000_M1 18000_30000_M1 0.020
r 18000_30000_M1 20000_30000_M1 0.020
r 20000_30000_M1 22000_30000_M1 0.020
r 22000_30000_M1 24000_30000_M1 0.020
r 24000_30000_M1 26000_30000_M1 0.020
r 26000_30000_M1 28000_30000_M1 0.020
r 28000_30000_M1 30000_30000_M1 0.020
r 30000_30000_M1 32000_30000_M1 0.020
r 32000_30000_M1 34000_30000_M1 0.020
r 34000_30000_M1 36000_30000_M1 0.020
r 36000_30000_M1 38000_30000_M1 0.020
r 38000_30000_M1 40000_30000_M1 0.020
r 40000_30000_M1 42000_30000_M1 0.020
r 42000_30000_M1 44000_30000_M1 0.020
r 44000_30000_M1 46000_30000_M1 0.020
r 46000_30000_M1 48000_30000_M1 0.020
r 48000_30000_M1 50000_30000_M1 0.020
r 50000_30000_M1 52000_30000_M1 0.020
r 52000_30000_M1 54000_30000_M1 0.020
r 54000_30000_M1 56000_30000_M1 0.020
r 56000_30000_M1 58000_30000_M1 0.020
r 58000_30000_M1 60000_30000_M1 0.020
r 60000_30000_M1 62000_30000_M1 0.020
r 62000_30000_M1 64000_30000_M1 0.020
r 64000_30000_M1 66000_30000_M1 0.020
r 66000_30000_M1 68000_30000_M1 0.020
r 68000_30000_M1 70000_30000_M1 0.020
r 70000_30000_M1 72000_30000_M1 0.020
r 72000_30000_M1 74000_30000_M1 0.020
r 74000_30000_M1 76000_30000_M1 0.020
r 76000_30000_M1 78000_30000_M1 0.020
r 78000_30000_M1 80000_30000_M1 0.020
r 80000_30000_M1 82000_30000_M1 0.020
r 82000_30000_M1 84000_30000_M1 0.020
r 84000_30000_M1 86000_30000_M1 0.020
r 86000_30000_M1 88000_30000_M1 0.020
r 88000_30000_M1 90000_30000_M1 0.020
r 90000_30000_M1 92000_30000_M1 0.020
r 92000_30000_M1 94000_30000_M1 0.020
r 94000_30000_M1 96000_30000_M1 0.020
r 96000_30000_M1 98000_30000_M1 0.020
r 98000_30000_M1 100000_30000_M1 0.020
r 2000_32000_M1 4000_32000_M1 0.020
r 4000_32000_M1 6000_32000_M1 0.020
r 6000_32000_M1 8000_32000_M1 0.020
r 8000_32000_M1 10000_32000_M1 0.020
r 10000_32000_M1 12000_32000_M1 0.020
r 12000_32000_M1 14000_32000_M1 0.020
r 14000_32000_M1 16000_32000_M1 0.020
r 16000_32000_M1 18000_32000_M1 0.020
r 18000_32000_M1 20000_32000_M1 0.020
r 20000_32000_M1 22000_32000_M1 0.020
r 22000_32000_M1 24000_32000_M1 0.020
r 24000_32000_M1 26000_32000_M1 0.020
r 26000_32000_M1 28000_32000_M1 0.020
r 28000_32000_M1 30000_32000_M1 0.020
r 30000_32000_M1 32000_32000_M1 0.020
r 32000_32000_M1 34000_32000_M1 0.020
r 34000_32000_M1 36000_32000_M1 0.020
r 36000_32000_M1 38000_32000_M1 0.020
r 38000_32000_M1 40000_32000_M1 0.020
r 40000_32000_M1 42000_32000_M1 0.020
r 42000_32000_M1 44000_32000_M1 0.020
r 44000_32000_M1 46000_32000_M1 0.020
r 46000_32000_M1 48000_32000_M1 0.020
r 48000_32000_M1 50000_32000_M1 0.020
r 50000_32000_M1 52000_32000_M1 0.020
r 52000_32000_M1 54000_32000_M1 0.020
r 54000_32000_M1 56000_32000_M1 0.020
r 56000_32000_M1 58000_32000_M1 0.020
r 58000_32000_M1 60000_32000_M1 0.020
r 60000_32000_M1 62000_32000_M1 0.020
r 62000_32000_M1 64000_32000_M1 0.020
r 64000_32000_M1 66000_32000_M1 0.020
r 66000_32000_M1 68000_32000_M1 0.020
r 68000_32000_M1 70000_32000_M1 0.020
r 70000_32000_M1 72000_32000_M1 0.020
r 72000_32000_M1 74000_32000_M1 0.020
r 74000_32000_M1 76000_32000_M1 0.020
r 76000_32000_M1 78000_32000_M1 0.020
r 78000_32000_M1 80000_32000_M1 0.020
r 80000_32000_M1 82000_32000_M1 0.020
r 82000_32000_M1 84000_32000_M1 0.020
r 84000_32000_M1 86000_32000_M1 0.020
r 86000_32000_M1 88000_32000_M1 0.020
r 88000_32000_M1 90000_32000_M1 0.020
r 90000_32000_M1 92000_32000_M1 0.020
r 92000_32000_M1 94000_32000_M1 0.020
r 94000_32000_M1 96000_32000_M1 0.020
r 96000_32000_M1 98000_32000_M1 0.020
r 98000_32000_M1 100000_32000_M1 0.020
r 2000_34000_M1 4000_34000_M1 0.020
r 4000_34000_M1 6000_34000_M1 0.020
r 6000_34000_M1 8000_34000_M1 0.020
r 8000_34000_M1 10000_34000_M1 0.020
r 10000_34000_M1 12000_34000_M1 0.020
r 12000_34000_M1 14000_34000_M1 0.020
r 14000_34000_M1 16000_34000_M1 0.020
r 16000_34000_M1 18000_34000_M1 0.020
r 18000_34000_M1 20000_34000_M1 0.020
r 20000_34000_M1 22000_34000_M1 0.020
r 22000_34000_M1 24000_34000_M1 0.020
r 24000_34000_M1 26000_34000_M1 0.020
r 26000_34000_M1 28000_34000_M1 0.020
r 28000_34000_M1 30000_34000_M1 0.020
r 30000_34000_M1 32000_34000_M1 0.020
r 32000_34000_M1 34000_34000_M1 0.020
r 34000_34000_M1 36000_34000_M1 0.020
r 36000_34000_M1 38000_34000_M1 0.020
r 38000_34000_M1 40000_34000_M1 0.020
r 40000_34000_M1 42000_34000_M1 0.020
r 42000_34000_M1 44000_34000_M1 0.020
r 44000_34000_M1 46000_34000_M1 0.020
r 46000_34000_M1 48000_34000_M1 0.020
r 48000_34000_M1 50000_34000_M1 0.020
r 50000_34000_M1 52000_34000_M1 0.020
r 52000_34000_M1 54000_34000_M1 0.020
r 54000_34000_M1 56000_34000_M1 0.020
r 56000_34000_M1 58000_34000_M1 0.020
r 58000_34000_M1 60000_34000_M1 0.020
r 60000_34000_M1 62000_34000_M1 0.020
r 62000_34000_M1 64000_34000_M1 0.020
r 64000_34000_M1 66000_34000_M1 0.020
r 66000_34000_M1 68000_34000_M1 0.020
r 68000_34000_M1 70000_34000_M1 0.020
r 70000_34000_M1 72000_34000_M1 0.020
r 72000_34000_M1 74000_34000_M1 0.020
r 74000_34000_M1 76000_34000_M1 0.020
r 76000_34000_M1 78000_34000_M1 0.020
r 78000_34000_M1 80000_34000_M1 0.020
r 80000_34000_M1 82000_34000_M1 0.020
r 82000_34000_M1 84000_34000_M1 0.020
r 84000_34000_M1 86000_34000_M1 0.020
r 86000_34000_M1 88000_34000_M1 0.020
r 88000_34000_M1 90000_34000_M1 0.020
r 90000_34000_M1 92000_34000_M1 0.020
r 92000_34000_M1 94000_34000_M1 0.020
r 94000_34000_M1 96000_34000_M1 0.020
r 96000_34000_M1 98000_34000_M1 0.020
r 98000_34000_M1 100000_34000_M1 0.020
r 2000_36000_M1 4000_36000_M1 0.020
r 4000_36000_M1 6000_36000_M1 0.020
r 6000_36000_M1 8000_36000_M1 0.020
r 8000_36000_M1 10000_36000_M1 0.020
r 10000_36000_M1 12000_36000_M1 0.020
r 12000_36000_M1 14000_36000_M1 0.020
r 14000_36000_M1 16000_36000_M1 0.020
r 16000_36000_M1 18000_36000_M1 0.020
r 18000_36000_M1 20000_36000_M1 0.020
r 20000_36000_M1 22000_36000_M1 0.020
r 22000_36000_M1 24000_36000_M1 0.020
r 24000_36000_M1 26000_36000_M1 0.020
r 26000_36000_M1 28000_36000_M1 0.020
r 28000_36000_M1 30000_36000_M1 0.020
r 30000_36000_M1 32000_36000_M1 0.020
r 32000_36000_M1 34000_36000_M1 0.020
r 34000_36000_M1 36000_36000_M1 0.020
r 36000_36000_M1 38000_36000_M1 0.020
r 38000_36000_M1 40000_36000_M1 0.020
r 40000_36000_M1 42000_36000_M1 0.020
r 42000_36000_M1 44000_36000_M1 0.020
r 44000_36000_M1 46000_36000_M1 0.020
r 46000_36000_M1 48000_36000_M1 0.020
r 48000_36000_M1 50000_36000_M1 0.020
r 50000_36000_M1 52000_36000_M1 0.020
r 52000_36000_M1 54000_36000_M1 0.020
r 54000_36000_M1 56000_36000_M1 0.020
r 56000_36000_M1 58000_36000_M1 0.020
r 58000_36000_M1 60000_36000_M1 0.020
r 60000_36000_M1 62000_36000_M1 0.020
r 62000_36000_M1 64000_36000_M1 0.020
r 64000_36000_M1 66000_36000_M1 0.020
r 66000_36000_M1 68000_36000_M1 0.020
r 68000_36000_M1 70000_36000_M1 0.020
r 70000_36000_M1 72000_36000_M1 0.020
r 72000_36000_M1 74000_36000_M1 0.020
r 74000_36000_M1 76000_36000_M1 0.020
r 76000_36000_M1 78000_36000_M1 0.020
r 78000_36000_M1 80000_36000_M1 0.020
r 80000_36000_M1 82000_36000_M1 0.020
r 82000_36000_M1 84000_36000_M1 0.020
r 84000_36000_M1 86000_36000_M1 0.020
r 86000_36000_M1 88000_36000_M1 0.020
r 88000_36000_M1 90000_36000_M1 0.020
r 90000_36000_M1 92000_36000_M1 0.020
r 92000_36000_M1 94000_36000_M1 0.020
r 94000_36000_M1 96000_36000_M1 0.020
r 96000_36000_M1 98000_36000_M1 0.020
r 98000_36000_M1 100000_36000_M1 0.020
r 2000_38000_M1 4000_38000_M1 0.020
r 4000_38000_M1 6000_38000_M1 0.020
r 6000_38000_M1 8000_38000_M1 0.020
r 8000_38000_M1 10000_38000_M1 0.020
r 10000_38000_M1 12000_38000_M1 0.020
r 12000_38000_M1 14000_38000_M1 0.020
r 14000_38000_M1 16000_38000_M1 0.020
r 16000_38000_M1 18000_38000_M1 0.020
r 18000_38000_M1 20000_38000_M1 0.020
r 20000_38000_M1 22000_38000_M1 0.020
r 22000_38000_M1 24000_38000_M1 0.020
r 24000_38000_M1 26000_38000_M1 0.020
r 26000_38000_M1 28000_38000_M1 0.020
r 28000_38000_M1 30000_38000_M1 0.020
r 30000_38000_M1 32000_38000_M1 0.020
r 32000_38000_M1 34000_38000_M1 0.020
r 34000_38000_M1 36000_38000_M1 0.020
r 36000_38000_M1 38000_38000_M1 0.020
r 38000_38000_M1 40000_38000_M1 0.020
r 40000_38000_M1 42000_38000_M1 0.020
r 42000_38000_M1 44000_38000_M1 0.020
r 44000_38000_M1 46000_38000_M1 0.020
r 46000_38000_M1 48000_38000_M1 0.020
r 48000_38000_M1 50000_38000_M1 0.020
r 50000_38000_M1 52000_38000_M1 0.020
r 52000_38000_M1 54000_38000_M1 0.020
r 54000_38000_M1 56000_38000_M1 0.020
r 56000_38000_M1 58000_38000_M1 0.020
r 58000_38000_M1 60000_38000_M1 0.020
r 60000_38000_M1 62000_38000_M1 0.020
r 62000_38000_M1 64000_38000_M1 0.020
r 64000_38000_M1 66000_38000_M1 0.020
r 66000_38000_M1 68000_38000_M1 0.020
r 68000_38000_M1 70000_38000_M1 0.020
r 70000_38000_M1 72000_38000_M1 0.020
r 72000_38000_M1 74000_38000_M1 0.020
r 74000_38000_M1 76000_38000_M1 0.020
r 76000_38000_M1 78000_38000_M1 0.020
r 78000_38000_M1 80000_38000_M1 0.020
r 80000_38000_M1 82000_38000_M1 0.020
r 82000_38000_M1 84000_38000_M1 0.020
r 84000_38000_M1 86000_38000_M1 0.020
r 86000_38000_M1 88000_38000_M1 0.020
r 88000_38000_M1 90000_38000_M1 0.020
r 90000_38000_M1 92000_38000_M1 0.020
r 92000_38000_M1 94000_38000_M1 0.020
r 94000_38000_M1 96000_38000_M1 0.020
r 96000_38000_M1 98000_38000_M1 0.020
r 98000_38000_M1 100000_38000_M1 0.020
r 2000_40000_M1 4000_40000_M1 0.020
r 4000_40000_M1 6000_40000_M1 0.020
r 6000_40000_M1 8000_40000_M1 0.020
r 8000_40000_M1 10000_40000_M1 0.020
r 10000_40000_M1 12000_40000_M1 0.020
r 12000_40000_M1 14000_40000_M1 0.020
r 14000_40000_M1 16000_40000_M1 0.020
r 16000_40000_M1 18000_40000_M1 0.020
r 18000_40000_M1 20000_40000_M1 0.020
r 20000_40000_M1 22000_40000_M1 0.020
r 22000_40000_M1 24000_40000_M1 0.020
r 24000_40000_M1 26000_40000_M1 0.020
r 26000_40000_M1 28000_40000_M1 0.020
r 28000_40000_M1 30000_40000_M1 0.020
r 30000_40000_M1 32000_40000_M1 0.020
r 32000_40000_M1 34000_40000_M1 0.020
r 34000_40000_M1 36000_40000_M1 0.020
r 36000_40000_M1 38000_40000_M1 0.020
r 38000_40000_M1 40000_40000_M1 0.020
r 40000_40000_M1 42000_40000_M1 0.020
r 42000_40000_M1 44000_40000_M1 0.020
r 44000_40000_M1 46000_40000_M1 0.020
r 46000_40000_M1 48000_40000_M1 0.020
r 48000_40000_M1 50000_40000_M1 0.020
r 50000_40000_M1 52000_40000_M1 0.020
r 52000_40000_M1 54000_40000_M1 0.020
r 54000_40000_M1 56000_40000_M1 0.020
r 56000_40000_M1 58000_40000_M1 0.020
r 58000_40000_M1 60000_40000_M1 0.020
r 60000_40000_M1 62000_40000_M1 0.020
r 62000_40000_M1 64000_40000_M1 0.020
r 64000_40000_M1 66000_40000_M1 0.020
r 66000_40000_M1 68000_40000_M1 0.020
r 68000_40000_M1 70000_40000_M1 0.020
r 70000_40000_M1 72000_40000_M1 0.020
r 72000_40000_M1 74000_40000_M1 0.020
r 74000_40000_M1 76000_40000_M1 0.020
r 76000_40000_M1 78000_40000_M1 0.020
r 78000_40000_M1 80000_40000_M1 0.020
r 80000_40000_M1 82000_40000_M1 0.020
r 82000_40000_M1 84000_40000_M1 0.020
r 84000_40000_M1 86000_40000_M1 0.020
r 86000_40000_M1 88000_40000_M1 0.020
r 88000_40000_M1 90000_40000_M1 0.020
r 90000_40000_M1 92000_40000_M1 0.020
r 92000_40000_M1 94000_40000_M1 0.020
r 94000_40000_M1 96000_40000_M1 0.020
r 96000_40000_M1 98000_40000_M1 0.020
r 98000_40000_M1 100000_40000_M1 0.020
r 2000_42000_M1 4000_42000_M1 0.020
r 4000_42000_M1 6000_42000_M1 0.020
r 6000_42000_M1 8000_42000_M1 0.020
r 8000_42000_M1 10000_42000_M1 0.020
r 10000_42000_M1 12000_42000_M1 0.020
r 12000_42000_M1 14000_42000_M1 0.020
r 14000_42000_M1 16000_42000_M1 0.020
r 16000_42000_M1 18000_42000_M1 0.020
r 18000_42000_M1 20000_42000_M1 0.020
r 20000_42000_M1 22000_42000_M1 0.020
r 22000_42000_M1 24000_42000_M1 0.020
r 24000_42000_M1 26000_42000_M1 0.020
r 26000_42000_M1 28000_42000_M1 0.020
r 28000_42000_M1 30000_42000_M1 0.020
r 30000_42000_M1 32000_42000_M1 0.020
r 32000_42000_M1 34000_42000_M1 0.020
r 34000_42000_M1 36000_42000_M1 0.020
r 36000_42000_M1 38000_42000_M1 0.020
r 38000_42000_M1 40000_42000_M1 0.020
r 40000_42000_M1 42000_42000_M1 0.020
r 42000_42000_M1 44000_42000_M1 0.020
r 44000_42000_M1 46000_42000_M1 0.020
r 46000_42000_M1 48000_42000_M1 0.020
r 48000_42000_M1 50000_42000_M1 0.020
r 50000_42000_M1 52000_42000_M1 0.020
r 52000_42000_M1 54000_42000_M1 0.020
r 54000_42000_M1 56000_42000_M1 0.020
r 56000_42000_M1 58000_42000_M1 0.020
r 58000_42000_M1 60000_42000_M1 0.020
r 60000_42000_M1 62000_42000_M1 0.020
r 62000_42000_M1 64000_42000_M1 0.020
r 64000_42000_M1 66000_42000_M1 0.020
r 66000_42000_M1 68000_42000_M1 0.020
r 68000_42000_M1 70000_42000_M1 0.020
r 70000_42000_M1 72000_42000_M1 0.020
r 72000_42000_M1 74000_42000_M1 0.020
r 74000_42000_M1 76000_42000_M1 0.020
r 76000_42000_M1 78000_42000_M1 0.020
r 78000_42000_M1 80000_42000_M1 0.020
r 80000_42000_M1 82000_42000_M1 0.020
r 82000_42000_M1 84000_42000_M1 0.020
r 84000_42000_M1 86000_42000_M1 0.020
r 86000_42000_M1 88000_42000_M1 0.020
r 88000_42000_M1 90000_42000_M1 0.020
r 90000_42000_M1 92000_42000_M1 0.020
r 92000_42000_M1 94000_42000_M1 0.020
r 94000_42000_M1 96000_42000_M1 0.020
r 96000_42000_M1 98000_42000_M1 0.020
r 98000_42000_M1 100000_42000_M1 0.020
r 2000_44000_M1 4000_44000_M1 0.020
r 4000_44000_M1 6000_44000_M1 0.020
r 6000_44000_M1 8000_44000_M1 0.020
r 8000_44000_M1 10000_44000_M1 0.020
r 10000_44000_M1 12000_44000_M1 0.020
r 12000_44000_M1 14000_44000_M1 0.020
r 14000_44000_M1 16000_44000_M1 0.020
r 16000_44000_M1 18000_44000_M1 0.020
r 18000_44000_M1 20000_44000_M1 0.020
r 20000_44000_M1 22000_44000_M1 0.020
r 22000_44000_M1 24000_44000_M1 0.020
r 24000_44000_M1 26000_44000_M1 0.020
r 26000_44000_M1 28000_44000_M1 0.020
r 28000_44000_M1 30000_44000_M1 0.020
r 30000_44000_M1 32000_44000_M1 0.020
r 32000_44000_M1 34000_44000_M1 0.020
r 34000_44000_M1 36000_44000_M1 0.020
r 36000_44000_M1 38000_44000_M1 0.020
r 38000_44000_M1 40000_44000_M1 0.020
r 40000_44000_M1 42000_44000_M1 0.020
r 42000_44000_M1 44000_44000_M1 0.020
r 44000_44000_M1 46000_44000_M1 0.020
r 46000_44000_M1 48000_44000_M1 0.020
r 48000_44000_M1 50000_44000_M1 0.020
r 50000_44000_M1 52000_44000_M1 0.020
r 52000_44000_M1 54000_44000_M1 0.020
r 54000_44000_M1 56000_44000_M1 0.020
r 56000_44000_M1 58000_44000_M1 0.020
r 58000_44000_M1 60000_44000_M1 0.020
r 60000_44000_M1 62000_44000_M1 0.020
r 62000_44000_M1 64000_44000_M1 0.020
r 64000_44000_M1 66000_44000_M1 0.020
r 66000_44000_M1 68000_44000_M1 0.020
r 68000_44000_M1 70000_44000_M1 0.020
r 70000_44000_M1 72000_44000_M1 0.020
r 72000_44000_M1 74000_44000_M1 0.020
r 74000_44000_M1 76000_44000_M1 0.020
r 76000_44000_M1 78000_44000_M1 0.020
r 78000_44000_M1 80000_44000_M1 0.020
r 80000_44000_M1 82000_44000_M1 0.020
r 82000_44000_M1 84000_44000_M1 0.020
r 84000_44000_M1 86000_44000_M1 0.020
r 86000_44000_M1 88000_44000_M1 0.020
r 88000_44000_M1 90000_44000_M1 0.020
r 90000_44000_M1 92000_44000_M1 0.020
r 92000_44000_M1 94000_44000_M1 0.020
r 94000_44000_M1 96000_44000_M1 0.020
r 96000_44000_M1 98000_44000_M1 0.020
r 98000_44000_M1 100000_44000_M1 0.020
r 2000_46000_M1 4000_46000_M1 0.020
r 4000_46000_M1 6000_46000_M1 0.020
r 6000_46000_M1 8000_46000_M1 0.020
r 8000_46000_M1 10000_46000_M1 0.020
r 10000_46000_M1 12000_46000_M1 0.020
r 12000_46000_M1 14000_46000_M1 0.020
r 14000_46000_M1 16000_46000_M1 0.020
r 16000_46000_M1 18000_46000_M1 0.020
r 18000_46000_M1 20000_46000_M1 0.020
r 20000_46000_M1 22000_46000_M1 0.020
r 22000_46000_M1 24000_46000_M1 0.020
r 24000_46000_M1 26000_46000_M1 0.020
r 26000_46000_M1 28000_46000_M1 0.020
r 28000_46000_M1 30000_46000_M1 0.020
r 30000_46000_M1 32000_46000_M1 0.020
r 32000_46000_M1 34000_46000_M1 0.020
r 34000_46000_M1 36000_46000_M1 0.020
r 36000_46000_M1 38000_46000_M1 0.020
r 38000_46000_M1 40000_46000_M1 0.020
r 40000_46000_M1 42000_46000_M1 0.020
r 42000_46000_M1 44000_46000_M1 0.020
r 44000_46000_M1 46000_46000_M1 0.020
r 46000_46000_M1 48000_46000_M1 0.020
r 48000_46000_M1 50000_46000_M1 0.020
r 50000_46000_M1 52000_46000_M1 0.020
r 52000_46000_M1 54000_46000_M1 0.020
r 54000_46000_M1 56000_46000_M1 0.020
r 56000_46000_M1 58000_46000_M1 0.020
r 58000_46000_M1 60000_46000_M1 0.020
r 60000_46000_M1 62000_46000_M1 0.020
r 62000_46000_M1 64000_46000_M1 0.020
r 64000_46000_M1 66000_46000_M1 0.020
r 66000_46000_M1 68000_46000_M1 0.020
r 68000_46000_M1 70000_46000_M1 0.020
r 70000_46000_M1 72000_46000_M1 0.020
r 72000_46000_M1 74000_46000_M1 0.020
r 74000_46000_M1 76000_46000_M1 0.020
r 76000_46000_M1 78000_46000_M1 0.020
r 78000_46000_M1 80000_46000_M1 0.020
r 80000_46000_M1 82000_46000_M1 0.020
r 82000_46000_M1 84000_46000_M1 0.020
r 84000_46000_M1 86000_46000_M1 0.020
r 86000_46000_M1 88000_46000_M1 0.020
r 88000_46000_M1 90000_46000_M1 0.020
r 90000_46000_M1 92000_46000_M1 0.020
r 92000_46000_M1 94000_46000_M1 0.020
r 94000_46000_M1 96000_46000_M1 0.020
r 96000_46000_M1 98000_46000_M1 0.020
r 98000_46000_M1 100000_46000_M1 0.020
r 2000_48000_M1 4000_48000_M1 0.020
r 4000_48000_M1 6000_48000_M1 0.020
r 6000_48000_M1 8000_48000_M1 0.020
r 8000_48000_M1 10000_48000_M1 0.020
r 10000_48000_M1 12000_48000_M1 0.020
r 12000_48000_M1 14000_48000_M1 0.020
r 14000_48000_M1 16000_48000_M1 0.020
r 16000_48000_M1 18000_48000_M1 0.020
r 18000_48000_M1 20000_48000_M1 0.020
r 20000_48000_M1 22000_48000_M1 0.020
r 22000_48000_M1 24000_48000_M1 0.020
r 24000_48000_M1 26000_48000_M1 0.020
r 26000_48000_M1 28000_48000_M1 0.020
r 28000_48000_M1 30000_48000_M1 0.020
r 30000_48000_M1 32000_48000_M1 0.020
r 32000_48000_M1 34000_48000_M1 0.020
r 34000_48000_M1 36000_48000_M1 0.020
r 36000_48000_M1 38000_48000_M1 0.020
r 38000_48000_M1 40000_48000_M1 0.020
r 40000_48000_M1 42000_48000_M1 0.020
r 42000_48000_M1 44000_48000_M1 0.020
r 44000_48000_M1 46000_48000_M1 0.020
r 46000_48000_M1 48000_48000_M1 0.020
r 48000_48000_M1 50000_48000_M1 0.020
r 50000_48000_M1 52000_48000_M1 0.020
r 52000_48000_M1 54000_48000_M1 0.020
r 54000_48000_M1 56000_48000_M1 0.020
r 56000_48000_M1 58000_48000_M1 0.020
r 58000_48000_M1 60000_48000_M1 0.020
r 60000_48000_M1 62000_48000_M1 0.020
r 62000_48000_M1 64000_48000_M1 0.020
r 64000_48000_M1 66000_48000_M1 0.020
r 66000_48000_M1 68000_48000_M1 0.020
r 68000_48000_M1 70000_48000_M1 0.020
r 70000_48000_M1 72000_48000_M1 0.020
r 72000_48000_M1 74000_48000_M1 0.020
r 74000_48000_M1 76000_48000_M1 0.020
r 76000_48000_M1 78000_48000_M1 0.020
r 78000_48000_M1 80000_48000_M1 0.020
r 80000_48000_M1 82000_48000_M1 0.020
r 82000_48000_M1 84000_48000_M1 0.020
r 84000_48000_M1 86000_48000_M1 0.020
r 86000_48000_M1 88000_48000_M1 0.020
r 88000_48000_M1 90000_48000_M1 0.020
r 90000_48000_M1 92000_48000_M1 0.020
r 92000_48000_M1 94000_48000_M1 0.020
r 94000_48000_M1 96000_48000_M1 0.020
r 96000_48000_M1 98000_48000_M1 0.020
r 98000_48000_M1 100000_48000_M1 0.020
r 2000_50000_M1 4000_50000_M1 0.020
r 4000_50000_M1 6000_50000_M1 0.020
r 6000_50000_M1 8000_50000_M1 0.020
r 8000_50000_M1 10000_50000_M1 0.020
r 10000_50000_M1 12000_50000_M1 0.020
r 12000_50000_M1 14000_50000_M1 0.020
r 14000_50000_M1 16000_50000_M1 0.020
r 16000_50000_M1 18000_50000_M1 0.020
r 18000_50000_M1 20000_50000_M1 0.020
r 20000_50000_M1 22000_50000_M1 0.020
r 22000_50000_M1 24000_50000_M1 0.020
r 24000_50000_M1 26000_50000_M1 0.020
r 26000_50000_M1 28000_50000_M1 0.020
r 28000_50000_M1 30000_50000_M1 0.020
r 30000_50000_M1 32000_50000_M1 0.020
r 32000_50000_M1 34000_50000_M1 0.020
r 34000_50000_M1 36000_50000_M1 0.020
r 36000_50000_M1 38000_50000_M1 0.020
r 38000_50000_M1 40000_50000_M1 0.020
r 40000_50000_M1 42000_50000_M1 0.020
r 42000_50000_M1 44000_50000_M1 0.020
r 44000_50000_M1 46000_50000_M1 0.020
r 46000_50000_M1 48000_50000_M1 0.020
r 48000_50000_M1 50000_50000_M1 0.020
r 50000_50000_M1 52000_50000_M1 0.020
r 52000_50000_M1 54000_50000_M1 0.020
r 54000_50000_M1 56000_50000_M1 0.020
r 56000_50000_M1 58000_50000_M1 0.020
r 58000_50000_M1 60000_50000_M1 0.020
r 60000_50000_M1 62000_50000_M1 0.020
r 62000_50000_M1 64000_50000_M1 0.020
r 64000_50000_M1 66000_50000_M1 0.020
r 66000_50000_M1 68000_50000_M1 0.020
r 68000_50000_M1 70000_50000_M1 0.020
r 70000_50000_M1 72000_50000_M1 0.020
r 72000_50000_M1 74000_50000_M1 0.020
r 74000_50000_M1 76000_50000_M1 0.020
r 76000_50000_M1 78000_50000_M1 0.020
r 78000_50000_M1 80000_50000_M1 0.020
r 80000_50000_M1 82000_50000_M1 0.020
r 82000_50000_M1 84000_50000_M1 0.020
r 84000_50000_M1 86000_50000_M1 0.020
r 86000_50000_M1 88000_50000_M1 0.020
r 88000_50000_M1 90000_50000_M1 0.020
r 90000_50000_M1 92000_50000_M1 0.020
r 92000_50000_M1 94000_50000_M1 0.020
r 94000_50000_M1 96000_50000_M1 0.020
r 96000_50000_M1 98000_50000_M1 0.020
r 98000_50000_M1 100000_50000_M1 0.020
r 2000_52000_M1 4000_52000_M1 0.020
r 4000_52000_M1 6000_52000_M1 0.020
r 6000_52000_M1 8000_52000_M1 0.020
r 8000_52000_M1 10000_52000_M1 0.020
r 10000_52000_M1 12000_52000_M1 0.020
r 12000_52000_M1 14000_52000_M1 0.020
r 14000_52000_M1 16000_52000_M1 0.020
r 16000_52000_M1 18000_52000_M1 0.020
r 18000_52000_M1 20000_52000_M1 0.020
r 20000_52000_M1 22000_52000_M1 0.020
r 22000_52000_M1 24000_52000_M1 0.020
r 24000_52000_M1 26000_52000_M1 0.020
r 26000_52000_M1 28000_52000_M1 0.020
r 28000_52000_M1 30000_52000_M1 0.020
r 30000_52000_M1 32000_52000_M1 0.020
r 32000_52000_M1 34000_52000_M1 0.020
r 34000_52000_M1 36000_52000_M1 0.020
r 36000_52000_M1 38000_52000_M1 0.020
r 38000_52000_M1 40000_52000_M1 0.020
r 40000_52000_M1 42000_52000_M1 0.020
r 42000_52000_M1 44000_52000_M1 0.020
r 44000_52000_M1 46000_52000_M1 0.020
r 46000_52000_M1 48000_52000_M1 0.020
r 48000_52000_M1 50000_52000_M1 0.020
r 50000_52000_M1 52000_52000_M1 0.020
r 52000_52000_M1 54000_52000_M1 0.020
r 54000_52000_M1 56000_52000_M1 0.020
r 56000_52000_M1 58000_52000_M1 0.020
r 58000_52000_M1 60000_52000_M1 0.020
r 60000_52000_M1 62000_52000_M1 0.020
r 62000_52000_M1 64000_52000_M1 0.020
r 64000_52000_M1 66000_52000_M1 0.020
r 66000_52000_M1 68000_52000_M1 0.020
r 68000_52000_M1 70000_52000_M1 0.020
r 70000_52000_M1 72000_52000_M1 0.020
r 72000_52000_M1 74000_52000_M1 0.020
r 74000_52000_M1 76000_52000_M1 0.020
r 76000_52000_M1 78000_52000_M1 0.020
r 78000_52000_M1 80000_52000_M1 0.020
r 80000_52000_M1 82000_52000_M1 0.020
r 82000_52000_M1 84000_52000_M1 0.020
r 84000_52000_M1 86000_52000_M1 0.020
r 86000_52000_M1 88000_52000_M1 0.020
r 88000_52000_M1 90000_52000_M1 0.020
r 90000_52000_M1 92000_52000_M1 0.020
r 92000_52000_M1 94000_52000_M1 0.020
r 94000_52000_M1 96000_52000_M1 0.020
r 96000_52000_M1 98000_52000_M1 0.020
r 98000_52000_M1 100000_52000_M1 0.020
r 2000_54000_M1 4000_54000_M1 0.020
r 4000_54000_M1 6000_54000_M1 0.020
r 6000_54000_M1 8000_54000_M1 0.020
r 8000_54000_M1 10000_54000_M1 0.020
r 10000_54000_M1 12000_54000_M1 0.020
r 12000_54000_M1 14000_54000_M1 0.020
r 14000_54000_M1 16000_54000_M1 0.020
r 16000_54000_M1 18000_54000_M1 0.020
r 18000_54000_M1 20000_54000_M1 0.020
r 20000_54000_M1 22000_54000_M1 0.020
r 22000_54000_M1 24000_54000_M1 0.020
r 24000_54000_M1 26000_54000_M1 0.020
r 26000_54000_M1 28000_54000_M1 0.020
r 28000_54000_M1 30000_54000_M1 0.020
r 30000_54000_M1 32000_54000_M1 0.020
r 32000_54000_M1 34000_54000_M1 0.020
r 34000_54000_M1 36000_54000_M1 0.020
r 36000_54000_M1 38000_54000_M1 0.020
r 38000_54000_M1 40000_54000_M1 0.020
r 40000_54000_M1 42000_54000_M1 0.020
r 42000_54000_M1 44000_54000_M1 0.020
r 44000_54000_M1 46000_54000_M1 0.020
r 46000_54000_M1 48000_54000_M1 0.020
r 48000_54000_M1 50000_54000_M1 0.020
r 50000_54000_M1 52000_54000_M1 0.020
r 52000_54000_M1 54000_54000_M1 0.020
r 54000_54000_M1 56000_54000_M1 0.020
r 56000_54000_M1 58000_54000_M1 0.020
r 58000_54000_M1 60000_54000_M1 0.020
r 60000_54000_M1 62000_54000_M1 0.020
r 62000_54000_M1 64000_54000_M1 0.020
r 64000_54000_M1 66000_54000_M1 0.020
r 66000_54000_M1 68000_54000_M1 0.020
r 68000_54000_M1 70000_54000_M1 0.020
r 70000_54000_M1 72000_54000_M1 0.020
r 72000_54000_M1 74000_54000_M1 0.020
r 74000_54000_M1 76000_54000_M1 0.020
r 76000_54000_M1 78000_54000_M1 0.020
r 78000_54000_M1 80000_54000_M1 0.020
r 80000_54000_M1 82000_54000_M1 0.020
r 82000_54000_M1 84000_54000_M1 0.020
r 84000_54000_M1 86000_54000_M1 0.020
r 86000_54000_M1 88000_54000_M1 0.020
r 88000_54000_M1 90000_54000_M1 0.020
r 90000_54000_M1 92000_54000_M1 0.020
r 92000_54000_M1 94000_54000_M1 0.020
r 94000_54000_M1 96000_54000_M1 0.020
r 96000_54000_M1 98000_54000_M1 0.020
r 98000_54000_M1 100000_54000_M1 0.020
r 2000_56000_M1 4000_56000_M1 0.020
r 4000_56000_M1 6000_56000_M1 0.020
r 6000_56000_M1 8000_56000_M1 0.020
r 8000_56000_M1 10000_56000_M1 0.020
r 10000_56000_M1 12000_56000_M1 0.020
r 12000_56000_M1 14000_56000_M1 0.020
r 14000_56000_M1 16000_56000_M1 0.020
r 16000_56000_M1 18000_56000_M1 0.020
r 18000_56000_M1 20000_56000_M1 0.020
r 20000_56000_M1 22000_56000_M1 0.020
r 22000_56000_M1 24000_56000_M1 0.020
r 24000_56000_M1 26000_56000_M1 0.020
r 26000_56000_M1 28000_56000_M1 0.020
r 28000_56000_M1 30000_56000_M1 0.020
r 30000_56000_M1 32000_56000_M1 0.020
r 32000_56000_M1 34000_56000_M1 0.020
r 34000_56000_M1 36000_56000_M1 0.020
r 36000_56000_M1 38000_56000_M1 0.020
r 38000_56000_M1 40000_56000_M1 0.020
r 40000_56000_M1 42000_56000_M1 0.020
r 42000_56000_M1 44000_56000_M1 0.020
r 44000_56000_M1 46000_56000_M1 0.020
r 46000_56000_M1 48000_56000_M1 0.020
r 48000_56000_M1 50000_56000_M1 0.020
r 50000_56000_M1 52000_56000_M1 0.020
r 52000_56000_M1 54000_56000_M1 0.020
r 54000_56000_M1 56000_56000_M1 0.020
r 56000_56000_M1 58000_56000_M1 0.020
r 58000_56000_M1 60000_56000_M1 0.020
r 60000_56000_M1 62000_56000_M1 0.020
r 62000_56000_M1 64000_56000_M1 0.020
r 64000_56000_M1 66000_56000_M1 0.020
r 66000_56000_M1 68000_56000_M1 0.020
r 68000_56000_M1 70000_56000_M1 0.020
r 70000_56000_M1 72000_56000_M1 0.020
r 72000_56000_M1 74000_56000_M1 0.020
r 74000_56000_M1 76000_56000_M1 0.020
r 76000_56000_M1 78000_56000_M1 0.020
r 78000_56000_M1 80000_56000_M1 0.020
r 80000_56000_M1 82000_56000_M1 0.020
r 82000_56000_M1 84000_56000_M1 0.020
r 84000_56000_M1 86000_56000_M1 0.020
r 86000_56000_M1 88000_56000_M1 0.020
r 88000_56000_M1 90000_56000_M1 0.020
r 90000_56000_M1 92000_56000_M1 0.020
r 92000_56000_M1 94000_56000_M1 0.020
r 94000_56000_M1 96000_56000_M1 0.020
r 96000_56000_M1 98000_56000_M1 0.020
r 98000_56000_M1 100000_56000_M1 0.020
r 2000_58000_M1 4000_58000_M1 0.020
r 4000_58000_M1 6000_58000_M1 0.020
r 6000_58000_M1 8000_58000_M1 0.020
r 8000_58000_M1 10000_58000_M1 0.020
r 10000_58000_M1 12000_58000_M1 0.020
r 12000_58000_M1 14000_58000_M1 0.020
r 14000_58000_M1 16000_58000_M1 0.020
r 16000_58000_M1 18000_58000_M1 0.020
r 18000_58000_M1 20000_58000_M1 0.020
r 20000_58000_M1 22000_58000_M1 0.020
r 22000_58000_M1 24000_58000_M1 0.020
r 24000_58000_M1 26000_58000_M1 0.020
r 26000_58000_M1 28000_58000_M1 0.020
r 28000_58000_M1 30000_58000_M1 0.020
r 30000_58000_M1 32000_58000_M1 0.020
r 32000_58000_M1 34000_58000_M1 0.020
r 34000_58000_M1 36000_58000_M1 0.020
r 36000_58000_M1 38000_58000_M1 0.020
r 38000_58000_M1 40000_58000_M1 0.020
r 40000_58000_M1 42000_58000_M1 0.020
r 42000_58000_M1 44000_58000_M1 0.020
r 44000_58000_M1 46000_58000_M1 0.020
r 46000_58000_M1 48000_58000_M1 0.020
r 48000_58000_M1 50000_58000_M1 0.020
r 50000_58000_M1 52000_58000_M1 0.020
r 52000_58000_M1 54000_58000_M1 0.020
r 54000_58000_M1 56000_58000_M1 0.020
r 56000_58000_M1 58000_58000_M1 0.020
r 58000_58000_M1 60000_58000_M1 0.020
r 60000_58000_M1 62000_58000_M1 0.020
r 62000_58000_M1 64000_58000_M1 0.020
r 64000_58000_M1 66000_58000_M1 0.020
r 66000_58000_M1 68000_58000_M1 0.020
r 68000_58000_M1 70000_58000_M1 0.020
r 70000_58000_M1 72000_58000_M1 0.020
r 72000_58000_M1 74000_58000_M1 0.020
r 74000_58000_M1 76000_58000_M1 0.020
r 76000_58000_M1 78000_58000_M1 0.020
r 78000_58000_M1 80000_58000_M1 0.020
r 80000_58000_M1 82000_58000_M1 0.020
r 82000_58000_M1 84000_58000_M1 0.020
r 84000_58000_M1 86000_58000_M1 0.020
r 86000_58000_M1 88000_58000_M1 0.020
r 88000_58000_M1 90000_58000_M1 0.020
r 90000_58000_M1 92000_58000_M1 0.020
r 92000_58000_M1 94000_58000_M1 0.020
r 94000_58000_M1 96000_58000_M1 0.020
r 96000_58000_M1 98000_58000_M1 0.020
r 98000_58000_M1 100000_58000_M1 0.020
r 2000_60000_M1 4000_60000_M1 0.020
r 4000_60000_M1 6000_60000_M1 0.020
r 6000_60000_M1 8000_60000_M1 0.020
r 8000_60000_M1 10000_60000_M1 0.020
r 10000_60000_M1 12000_60000_M1 0.020
r 12000_60000_M1 14000_60000_M1 0.020
r 14000_60000_M1 16000_60000_M1 0.020
r 16000_60000_M1 18000_60000_M1 0.020
r 18000_60000_M1 20000_60000_M1 0.020
r 20000_60000_M1 22000_60000_M1 0.020
r 22000_60000_M1 24000_60000_M1 0.020
r 24000_60000_M1 26000_60000_M1 0.020
r 26000_60000_M1 28000_60000_M1 0.020
r 28000_60000_M1 30000_60000_M1 0.020
r 30000_60000_M1 32000_60000_M1 0.020
r 32000_60000_M1 34000_60000_M1 0.020
r 34000_60000_M1 36000_60000_M1 0.020
r 36000_60000_M1 38000_60000_M1 0.020
r 38000_60000_M1 40000_60000_M1 0.020
r 40000_60000_M1 42000_60000_M1 0.020
r 42000_60000_M1 44000_60000_M1 0.020
r 44000_60000_M1 46000_60000_M1 0.020
r 46000_60000_M1 48000_60000_M1 0.020
r 48000_60000_M1 50000_60000_M1 0.020
r 50000_60000_M1 52000_60000_M1 0.020
r 52000_60000_M1 54000_60000_M1 0.020
r 54000_60000_M1 56000_60000_M1 0.020
r 56000_60000_M1 58000_60000_M1 0.020
r 58000_60000_M1 60000_60000_M1 0.020
r 60000_60000_M1 62000_60000_M1 0.020
r 62000_60000_M1 64000_60000_M1 0.020
r 64000_60000_M1 66000_60000_M1 0.020
r 66000_60000_M1 68000_60000_M1 0.020
r 68000_60000_M1 70000_60000_M1 0.020
r 70000_60000_M1 72000_60000_M1 0.020
r 72000_60000_M1 74000_60000_M1 0.020
r 74000_60000_M1 76000_60000_M1 0.020
r 76000_60000_M1 78000_60000_M1 0.020
r 78000_60000_M1 80000_60000_M1 0.020
r 80000_60000_M1 82000_60000_M1 0.020
r 82000_60000_M1 84000_60000_M1 0.020
r 84000_60000_M1 86000_60000_M1 0.020
r 86000_60000_M1 88000_60000_M1 0.020
r 88000_60000_M1 90000_60000_M1 0.020
r 90000_60000_M1 92000_60000_M1 0.020
r 92000_60000_M1 94000_60000_M1 0.020
r 94000_60000_M1 96000_60000_M1 0.020
r 96000_60000_M1 98000_60000_M1 0.020
r 98000_60000_M1 100000_60000_M1 0.020
r 2000_62000_M1 4000_62000_M1 0.020
r 4000_62000_M1 6000_62000_M1 0.020
r 6000_62000_M1 8000_62000_M1 0.020
r 8000_62000_M1 10000_62000_M1 0.020
r 10000_62000_M1 12000_62000_M1 0.020
r 12000_62000_M1 14000_62000_M1 0.020
r 14000_62000_M1 16000_62000_M1 0.020
r 16000_62000_M1 18000_62000_M1 0.020
r 18000_62000_M1 20000_62000_M1 0.020
r 20000_62000_M1 22000_62000_M1 0.020
r 22000_62000_M1 24000_62000_M1 0.020
r 24000_62000_M1 26000_62000_M1 0.020
r 26000_62000_M1 28000_62000_M1 0.020
r 28000_62000_M1 30000_62000_M1 0.020
r 30000_62000_M1 32000_62000_M1 0.020
r 32000_62000_M1 34000_62000_M1 0.020
r 34000_62000_M1 36000_62000_M1 0.020
r 36000_62000_M1 38000_62000_M1 0.020
r 38000_62000_M1 40000_62000_M1 0.020
r 40000_62000_M1 42000_62000_M1 0.020
r 42000_62000_M1 44000_62000_M1 0.020
r 44000_62000_M1 46000_62000_M1 0.020
r 46000_62000_M1 48000_62000_M1 0.020
r 48000_62000_M1 50000_62000_M1 0.020
r 50000_62000_M1 52000_62000_M1 0.020
r 52000_62000_M1 54000_62000_M1 0.020
r 54000_62000_M1 56000_62000_M1 0.020
r 56000_62000_M1 58000_62000_M1 0.020
r 58000_62000_M1 60000_62000_M1 0.020
r 60000_62000_M1 62000_62000_M1 0.020
r 62000_62000_M1 64000_62000_M1 0.020
r 64000_62000_M1 66000_62000_M1 0.020
r 66000_62000_M1 68000_62000_M1 0.020
r 68000_62000_M1 70000_62000_M1 0.020
r 70000_62000_M1 72000_62000_M1 0.020
r 72000_62000_M1 74000_62000_M1 0.020
r 74000_62000_M1 76000_62000_M1 0.020
r 76000_62000_M1 78000_62000_M1 0.020
r 78000_62000_M1 80000_62000_M1 0.020
r 80000_62000_M1 82000_62000_M1 0.020
r 82000_62000_M1 84000_62000_M1 0.020
r 84000_62000_M1 86000_62000_M1 0.020
r 86000_62000_M1 88000_62000_M1 0.020
r 88000_62000_M1 90000_62000_M1 0.020
r 90000_62000_M1 92000_62000_M1 0.020
r 92000_62000_M1 94000_62000_M1 0.020
r 94000_62000_M1 96000_62000_M1 0.020
r 96000_62000_M1 98000_62000_M1 0.020
r 98000_62000_M1 100000_62000_M1 0.020
r 2000_64000_M1 4000_64000_M1 0.020
r 4000_64000_M1 6000_64000_M1 0.020
r 6000_64000_M1 8000_64000_M1 0.020
r 8000_64000_M1 10000_64000_M1 0.020
r 10000_64000_M1 12000_64000_M1 0.020
r 12000_64000_M1 14000_64000_M1 0.020
r 14000_64000_M1 16000_64000_M1 0.020
r 16000_64000_M1 18000_64000_M1 0.020
r 18000_64000_M1 20000_64000_M1 0.020
r 20000_64000_M1 22000_64000_M1 0.020
r 22000_64000_M1 24000_64000_M1 0.020
r 24000_64000_M1 26000_64000_M1 0.020
r 26000_64000_M1 28000_64000_M1 0.020
r 28000_64000_M1 30000_64000_M1 0.020
r 30000_64000_M1 32000_64000_M1 0.020
r 32000_64000_M1 34000_64000_M1 0.020
r 34000_64000_M1 36000_64000_M1 0.020
r 36000_64000_M1 38000_64000_M1 0.020
r 38000_64000_M1 40000_64000_M1 0.020
r 40000_64000_M1 42000_64000_M1 0.020
r 42000_64000_M1 44000_64000_M1 0.020
r 44000_64000_M1 46000_64000_M1 0.020
r 46000_64000_M1 48000_64000_M1 0.020
r 48000_64000_M1 50000_64000_M1 0.020
r 50000_64000_M1 52000_64000_M1 0.020
r 52000_64000_M1 54000_64000_M1 0.020
r 54000_64000_M1 56000_64000_M1 0.020
r 56000_64000_M1 58000_64000_M1 0.020
r 58000_64000_M1 60000_64000_M1 0.020
r 60000_64000_M1 62000_64000_M1 0.020
r 62000_64000_M1 64000_64000_M1 0.020
r 64000_64000_M1 66000_64000_M1 0.020
r 66000_64000_M1 68000_64000_M1 0.020
r 68000_64000_M1 70000_64000_M1 0.020
r 70000_64000_M1 72000_64000_M1 0.020
r 72000_64000_M1 74000_64000_M1 0.020
r 74000_64000_M1 76000_64000_M1 0.020
r 76000_64000_M1 78000_64000_M1 0.020
r 78000_64000_M1 80000_64000_M1 0.020
r 80000_64000_M1 82000_64000_M1 0.020
r 82000_64000_M1 84000_64000_M1 0.020
r 84000_64000_M1 86000_64000_M1 0.020
r 86000_64000_M1 88000_64000_M1 0.020
r 88000_64000_M1 90000_64000_M1 0.020
r 90000_64000_M1 92000_64000_M1 0.020
r 92000_64000_M1 94000_64000_M1 0.020
r 94000_64000_M1 96000_64000_M1 0.020
r 96000_64000_M1 98000_64000_M1 0.020
r 98000_64000_M1 100000_64000_M1 0.020
r 2000_66000_M1 4000_66000_M1 0.020
r 4000_66000_M1 6000_66000_M1 0.020
r 6000_66000_M1 8000_66000_M1 0.020
r 8000_66000_M1 10000_66000_M1 0.020
r 10000_66000_M1 12000_66000_M1 0.020
r 12000_66000_M1 14000_66000_M1 0.020
r 14000_66000_M1 16000_66000_M1 0.020
r 16000_66000_M1 18000_66000_M1 0.020
r 18000_66000_M1 20000_66000_M1 0.020
r 20000_66000_M1 22000_66000_M1 0.020
r 22000_66000_M1 24000_66000_M1 0.020
r 24000_66000_M1 26000_66000_M1 0.020
r 26000_66000_M1 28000_66000_M1 0.020
r 28000_66000_M1 30000_66000_M1 0.020
r 30000_66000_M1 32000_66000_M1 0.020
r 32000_66000_M1 34000_66000_M1 0.020
r 34000_66000_M1 36000_66000_M1 0.020
r 36000_66000_M1 38000_66000_M1 0.020
r 38000_66000_M1 40000_66000_M1 0.020
r 40000_66000_M1 42000_66000_M1 0.020
r 42000_66000_M1 44000_66000_M1 0.020
r 44000_66000_M1 46000_66000_M1 0.020
r 46000_66000_M1 48000_66000_M1 0.020
r 48000_66000_M1 50000_66000_M1 0.020
r 50000_66000_M1 52000_66000_M1 0.020
r 52000_66000_M1 54000_66000_M1 0.020
r 54000_66000_M1 56000_66000_M1 0.020
r 56000_66000_M1 58000_66000_M1 0.020
r 58000_66000_M1 60000_66000_M1 0.020
r 60000_66000_M1 62000_66000_M1 0.020
r 62000_66000_M1 64000_66000_M1 0.020
r 64000_66000_M1 66000_66000_M1 0.020
r 66000_66000_M1 68000_66000_M1 0.020
r 68000_66000_M1 70000_66000_M1 0.020
r 70000_66000_M1 72000_66000_M1 0.020
r 72000_66000_M1 74000_66000_M1 0.020
r 74000_66000_M1 76000_66000_M1 0.020
r 76000_66000_M1 78000_66000_M1 0.020
r 78000_66000_M1 80000_66000_M1 0.020
r 80000_66000_M1 82000_66000_M1 0.020
r 82000_66000_M1 84000_66000_M1 0.020
r 84000_66000_M1 86000_66000_M1 0.020
r 86000_66000_M1 88000_66000_M1 0.020
r 88000_66000_M1 90000_66000_M1 0.020
r 90000_66000_M1 92000_66000_M1 0.020
r 92000_66000_M1 94000_66000_M1 0.020
r 94000_66000_M1 96000_66000_M1 0.020
r 96000_66000_M1 98000_66000_M1 0.020
r 98000_66000_M1 100000_66000_M1 0.020
r 2000_68000_M1 4000_68000_M1 0.020
r 4000_68000_M1 6000_68000_M1 0.020
r 6000_68000_M1 8000_68000_M1 0.020
r 8000_68000_M1 10000_68000_M1 0.020
r 10000_68000_M1 12000_68000_M1 0.020
r 12000_68000_M1 14000_68000_M1 0.020
r 14000_68000_M1 16000_68000_M1 0.020
r 16000_68000_M1 18000_68000_M1 0.020
r 18000_68000_M1 20000_68000_M1 0.020
r 20000_68000_M1 22000_68000_M1 0.020
r 22000_68000_M1 24000_68000_M1 0.020
r 24000_68000_M1 26000_68000_M1 0.020
r 26000_68000_M1 28000_68000_M1 0.020
r 28000_68000_M1 30000_68000_M1 0.020
r 30000_68000_M1 32000_68000_M1 0.020
r 32000_68000_M1 34000_68000_M1 0.020
r 34000_68000_M1 36000_68000_M1 0.020
r 36000_68000_M1 38000_68000_M1 0.020
r 38000_68000_M1 40000_68000_M1 0.020
r 40000_68000_M1 42000_68000_M1 0.020
r 42000_68000_M1 44000_68000_M1 0.020
r 44000_68000_M1 46000_68000_M1 0.020
r 46000_68000_M1 48000_68000_M1 0.020
r 48000_68000_M1 50000_68000_M1 0.020
r 50000_68000_M1 52000_68000_M1 0.020
r 52000_68000_M1 54000_68000_M1 0.020
r 54000_68000_M1 56000_68000_M1 0.020
r 56000_68000_M1 58000_68000_M1 0.020
r 58000_68000_M1 60000_68000_M1 0.020
r 60000_68000_M1 62000_68000_M1 0.020
r 62000_68000_M1 64000_68000_M1 0.020
r 64000_68000_M1 66000_68000_M1 0.020
r 66000_68000_M1 68000_68000_M1 0.020
r 68000_68000_M1 70000_68000_M1 0.020
r 70000_68000_M1 72000_68000_M1 0.020
r 72000_68000_M1 74000_68000_M1 0.020
r 74000_68000_M1 76000_68000_M1 0.020
r 76000_68000_M1 78000_68000_M1 0.020
r 78000_68000_M1 80000_68000_M1 0.020
r 80000_68000_M1 82000_68000_M1 0.020
r 82000_68000_M1 84000_68000_M1 0.020
r 84000_68000_M1 86000_68000_M1 0.020
r 86000_68000_M1 88000_68000_M1 0.020
r 88000_68000_M1 90000_68000_M1 0.020
r 90000_68000_M1 92000_68000_M1 0.020
r 92000_68000_M1 94000_68000_M1 0.020
r 94000_68000_M1 96000_68000_M1 0.020
r 96000_68000_M1 98000_68000_M1 0.020
r 98000_68000_M1 100000_68000_M1 0.020
r 2000_70000_M1 4000_70000_M1 0.020
r 4000_70000_M1 6000_70000_M1 0.020
r 6000_70000_M1 8000_70000_M1 0.020
r 8000_70000_M1 10000_70000_M1 0.020
r 10000_70000_M1 12000_70000_M1 0.020
r 12000_70000_M1 14000_70000_M1 0.020
r 14000_70000_M1 16000_70000_M1 0.020
r 16000_70000_M1 18000_70000_M1 0.020
r 18000_70000_M1 20000_70000_M1 0.020
r 20000_70000_M1 22000_70000_M1 0.020
r 22000_70000_M1 24000_70000_M1 0.020
r 24000_70000_M1 26000_70000_M1 0.020
r 26000_70000_M1 28000_70000_M1 0.020
r 28000_70000_M1 30000_70000_M1 0.020
r 30000_70000_M1 32000_70000_M1 0.020
r 32000_70000_M1 34000_70000_M1 0.020
r 34000_70000_M1 36000_70000_M1 0.020
r 36000_70000_M1 38000_70000_M1 0.020
r 38000_70000_M1 40000_70000_M1 0.020
r 40000_70000_M1 42000_70000_M1 0.020
r 42000_70000_M1 44000_70000_M1 0.020
r 44000_70000_M1 46000_70000_M1 0.020
r 46000_70000_M1 48000_70000_M1 0.020
r 48000_70000_M1 50000_70000_M1 0.020
r 50000_70000_M1 52000_70000_M1 0.020
r 52000_70000_M1 54000_70000_M1 0.020
r 54000_70000_M1 56000_70000_M1 0.020
r 56000_70000_M1 58000_70000_M1 0.020
r 58000_70000_M1 60000_70000_M1 0.020
r 60000_70000_M1 62000_70000_M1 0.020
r 62000_70000_M1 64000_70000_M1 0.020
r 64000_70000_M1 66000_70000_M1 0.020
r 66000_70000_M1 68000_70000_M1 0.020
r 68000_70000_M1 70000_70000_M1 0.020
r 70000_70000_M1 72000_70000_M1 0.020
r 72000_70000_M1 74000_70000_M1 0.020
r 74000_70000_M1 76000_70000_M1 0.020
r 76000_70000_M1 78000_70000_M1 0.020
r 78000_70000_M1 80000_70000_M1 0.020
r 80000_70000_M1 82000_70000_M1 0.020
r 82000_70000_M1 84000_70000_M1 0.020
r 84000_70000_M1 86000_70000_M1 0.020
r 86000_70000_M1 88000_70000_M1 0.020
r 88000_70000_M1 90000_70000_M1 0.020
r 90000_70000_M1 92000_70000_M1 0.020
r 92000_70000_M1 94000_70000_M1 0.020
r 94000_70000_M1 96000_70000_M1 0.020
r 96000_70000_M1 98000_70000_M1 0.020
r 98000_70000_M1 100000_70000_M1 0.020
r 2000_72000_M1 4000_72000_M1 0.020
r 4000_72000_M1 6000_72000_M1 0.020
r 6000_72000_M1 8000_72000_M1 0.020
r 8000_72000_M1 10000_72000_M1 0.020
r 10000_72000_M1 12000_72000_M1 0.020
r 12000_72000_M1 14000_72000_M1 0.020
r 14000_72000_M1 16000_72000_M1 0.020
r 16000_72000_M1 18000_72000_M1 0.020
r 18000_72000_M1 20000_72000_M1 0.020
r 20000_72000_M1 22000_72000_M1 0.020
r 22000_72000_M1 24000_72000_M1 0.020
r 24000_72000_M1 26000_72000_M1 0.020
r 26000_72000_M1 28000_72000_M1 0.020
r 28000_72000_M1 30000_72000_M1 0.020
r 30000_72000_M1 32000_72000_M1 0.020
r 32000_72000_M1 34000_72000_M1 0.020
r 34000_72000_M1 36000_72000_M1 0.020
r 36000_72000_M1 38000_72000_M1 0.020
r 38000_72000_M1 40000_72000_M1 0.020
r 40000_72000_M1 42000_72000_M1 0.020
r 42000_72000_M1 44000_72000_M1 0.020
r 44000_72000_M1 46000_72000_M1 0.020
r 46000_72000_M1 48000_72000_M1 0.020
r 48000_72000_M1 50000_72000_M1 0.020
r 50000_72000_M1 52000_72000_M1 0.020
r 52000_72000_M1 54000_72000_M1 0.020
r 54000_72000_M1 56000_72000_M1 0.020
r 56000_72000_M1 58000_72000_M1 0.020
r 58000_72000_M1 60000_72000_M1 0.020
r 60000_72000_M1 62000_72000_M1 0.020
r 62000_72000_M1 64000_72000_M1 0.020
r 64000_72000_M1 66000_72000_M1 0.020
r 66000_72000_M1 68000_72000_M1 0.020
r 68000_72000_M1 70000_72000_M1 0.020
r 70000_72000_M1 72000_72000_M1 0.020
r 72000_72000_M1 74000_72000_M1 0.020
r 74000_72000_M1 76000_72000_M1 0.020
r 76000_72000_M1 78000_72000_M1 0.020
r 78000_72000_M1 80000_72000_M1 0.020
r 80000_72000_M1 82000_72000_M1 0.020
r 82000_72000_M1 84000_72000_M1 0.020
r 84000_72000_M1 86000_72000_M1 0.020
r 86000_72000_M1 88000_72000_M1 0.020
r 88000_72000_M1 90000_72000_M1 0.020
r 90000_72000_M1 92000_72000_M1 0.020
r 92000_72000_M1 94000_72000_M1 0.020
r 94000_72000_M1 96000_72000_M1 0.020
r 96000_72000_M1 98000_72000_M1 0.020
r 98000_72000_M1 100000_72000_M1 0.020
r 2000_74000_M1 4000_74000_M1 0.020
r 4000_74000_M1 6000_74000_M1 0.020
r 6000_74000_M1 8000_74000_M1 0.020
r 8000_74000_M1 10000_74000_M1 0.020
r 10000_74000_M1 12000_74000_M1 0.020
r 12000_74000_M1 14000_74000_M1 0.020
r 14000_74000_M1 16000_74000_M1 0.020
r 16000_74000_M1 18000_74000_M1 0.020
r 18000_74000_M1 20000_74000_M1 0.020
r 20000_74000_M1 22000_74000_M1 0.020
r 22000_74000_M1 24000_74000_M1 0.020
r 24000_74000_M1 26000_74000_M1 0.020
r 26000_74000_M1 28000_74000_M1 0.020
r 28000_74000_M1 30000_74000_M1 0.020
r 30000_74000_M1 32000_74000_M1 0.020
r 32000_74000_M1 34000_74000_M1 0.020
r 34000_74000_M1 36000_74000_M1 0.020
r 36000_74000_M1 38000_74000_M1 0.020
r 38000_74000_M1 40000_74000_M1 0.020
r 40000_74000_M1 42000_74000_M1 0.020
r 42000_74000_M1 44000_74000_M1 0.020
r 44000_74000_M1 46000_74000_M1 0.020
r 46000_74000_M1 48000_74000_M1 0.020
r 48000_74000_M1 50000_74000_M1 0.020
r 50000_74000_M1 52000_74000_M1 0.020
r 52000_74000_M1 54000_74000_M1 0.020
r 54000_74000_M1 56000_74000_M1 0.020
r 56000_74000_M1 58000_74000_M1 0.020
r 58000_74000_M1 60000_74000_M1 0.020
r 60000_74000_M1 62000_74000_M1 0.020
r 62000_74000_M1 64000_74000_M1 0.020
r 64000_74000_M1 66000_74000_M1 0.020
r 66000_74000_M1 68000_74000_M1 0.020
r 68000_74000_M1 70000_74000_M1 0.020
r 70000_74000_M1 72000_74000_M1 0.020
r 72000_74000_M1 74000_74000_M1 0.020
r 74000_74000_M1 76000_74000_M1 0.020
r 76000_74000_M1 78000_74000_M1 0.020
r 78000_74000_M1 80000_74000_M1 0.020
r 80000_74000_M1 82000_74000_M1 0.020
r 82000_74000_M1 84000_74000_M1 0.020
r 84000_74000_M1 86000_74000_M1 0.020
r 86000_74000_M1 88000_74000_M1 0.020
r 88000_74000_M1 90000_74000_M1 0.020
r 90000_74000_M1 92000_74000_M1 0.020
r 92000_74000_M1 94000_74000_M1 0.020
r 94000_74000_M1 96000_74000_M1 0.020
r 96000_74000_M1 98000_74000_M1 0.020
r 98000_74000_M1 100000_74000_M1 0.020
r 2000_76000_M1 4000_76000_M1 0.020
r 4000_76000_M1 6000_76000_M1 0.020
r 6000_76000_M1 8000_76000_M1 0.020
r 8000_76000_M1 10000_76000_M1 0.020
r 10000_76000_M1 12000_76000_M1 0.020
r 12000_76000_M1 14000_76000_M1 0.020
r 14000_76000_M1 16000_76000_M1 0.020
r 16000_76000_M1 18000_76000_M1 0.020
r 18000_76000_M1 20000_76000_M1 0.020
r 20000_76000_M1 22000_76000_M1 0.020
r 22000_76000_M1 24000_76000_M1 0.020
r 24000_76000_M1 26000_76000_M1 0.020
r 26000_76000_M1 28000_76000_M1 0.020
r 28000_76000_M1 30000_76000_M1 0.020
r 30000_76000_M1 32000_76000_M1 0.020
r 32000_76000_M1 34000_76000_M1 0.020
r 34000_76000_M1 36000_76000_M1 0.020
r 36000_76000_M1 38000_76000_M1 0.020
r 38000_76000_M1 40000_76000_M1 0.020
r 40000_76000_M1 42000_76000_M1 0.020
r 42000_76000_M1 44000_76000_M1 0.020
r 44000_76000_M1 46000_76000_M1 0.020
r 46000_76000_M1 48000_76000_M1 0.020
r 48000_76000_M1 50000_76000_M1 0.020
r 50000_76000_M1 52000_76000_M1 0.020
r 52000_76000_M1 54000_76000_M1 0.020
r 54000_76000_M1 56000_76000_M1 0.020
r 56000_76000_M1 58000_76000_M1 0.020
r 58000_76000_M1 60000_76000_M1 0.020
r 60000_76000_M1 62000_76000_M1 0.020
r 62000_76000_M1 64000_76000_M1 0.020
r 64000_76000_M1 66000_76000_M1 0.020
r 66000_76000_M1 68000_76000_M1 0.020
r 68000_76000_M1 70000_76000_M1 0.020
r 70000_76000_M1 72000_76000_M1 0.020
r 72000_76000_M1 74000_76000_M1 0.020
r 74000_76000_M1 76000_76000_M1 0.020
r 76000_76000_M1 78000_76000_M1 0.020
r 78000_76000_M1 80000_76000_M1 0.020
r 80000_76000_M1 82000_76000_M1 0.020
r 82000_76000_M1 84000_76000_M1 0.020
r 84000_76000_M1 86000_76000_M1 0.020
r 86000_76000_M1 88000_76000_M1 0.020
r 88000_76000_M1 90000_76000_M1 0.020
r 90000_76000_M1 92000_76000_M1 0.020
r 92000_76000_M1 94000_76000_M1 0.020
r 94000_76000_M1 96000_76000_M1 0.020
r 96000_76000_M1 98000_76000_M1 0.020
r 98000_76000_M1 100000_76000_M1 0.020
r 2000_78000_M1 4000_78000_M1 0.020
r 4000_78000_M1 6000_78000_M1 0.020
r 6000_78000_M1 8000_78000_M1 0.020
r 8000_78000_M1 10000_78000_M1 0.020
r 10000_78000_M1 12000_78000_M1 0.020
r 12000_78000_M1 14000_78000_M1 0.020
r 14000_78000_M1 16000_78000_M1 0.020
r 16000_78000_M1 18000_78000_M1 0.020
r 18000_78000_M1 20000_78000_M1 0.020
r 20000_78000_M1 22000_78000_M1 0.020
r 22000_78000_M1 24000_78000_M1 0.020
r 24000_78000_M1 26000_78000_M1 0.020
r 26000_78000_M1 28000_78000_M1 0.020
r 28000_78000_M1 30000_78000_M1 0.020
r 30000_78000_M1 32000_78000_M1 0.020
r 32000_78000_M1 34000_78000_M1 0.020
r 34000_78000_M1 36000_78000_M1 0.020
r 36000_78000_M1 38000_78000_M1 0.020
r 38000_78000_M1 40000_78000_M1 0.020
r 40000_78000_M1 42000_78000_M1 0.020
r 42000_78000_M1 44000_78000_M1 0.020
r 44000_78000_M1 46000_78000_M1 0.020
r 46000_78000_M1 48000_78000_M1 0.020
r 48000_78000_M1 50000_78000_M1 0.020
r 50000_78000_M1 52000_78000_M1 0.020
r 52000_78000_M1 54000_78000_M1 0.020
r 54000_78000_M1 56000_78000_M1 0.020
r 56000_78000_M1 58000_78000_M1 0.020
r 58000_78000_M1 60000_78000_M1 0.020
r 60000_78000_M1 62000_78000_M1 0.020
r 62000_78000_M1 64000_78000_M1 0.020
r 64000_78000_M1 66000_78000_M1 0.020
r 66000_78000_M1 68000_78000_M1 0.020
r 68000_78000_M1 70000_78000_M1 0.020
r 70000_78000_M1 72000_78000_M1 0.020
r 72000_78000_M1 74000_78000_M1 0.020
r 74000_78000_M1 76000_78000_M1 0.020
r 76000_78000_M1 78000_78000_M1 0.020
r 78000_78000_M1 80000_78000_M1 0.020
r 80000_78000_M1 82000_78000_M1 0.020
r 82000_78000_M1 84000_78000_M1 0.020
r 84000_78000_M1 86000_78000_M1 0.020
r 86000_78000_M1 88000_78000_M1 0.020
r 88000_78000_M1 90000_78000_M1 0.020
r 90000_78000_M1 92000_78000_M1 0.020
r 92000_78000_M1 94000_78000_M1 0.020
r 94000_78000_M1 96000_78000_M1 0.020
r 96000_78000_M1 98000_78000_M1 0.020
r 98000_78000_M1 100000_78000_M1 0.020
r 2000_80000_M1 4000_80000_M1 0.020
r 4000_80000_M1 6000_80000_M1 0.020
r 6000_80000_M1 8000_80000_M1 0.020
r 8000_80000_M1 10000_80000_M1 0.020
r 10000_80000_M1 12000_80000_M1 0.020
r 12000_80000_M1 14000_80000_M1 0.020
r 14000_80000_M1 16000_80000_M1 0.020
r 16000_80000_M1 18000_80000_M1 0.020
r 18000_80000_M1 20000_80000_M1 0.020
r 20000_80000_M1 22000_80000_M1 0.020
r 22000_80000_M1 24000_80000_M1 0.020
r 24000_80000_M1 26000_80000_M1 0.020
r 26000_80000_M1 28000_80000_M1 0.020
r 28000_80000_M1 30000_80000_M1 0.020
r 30000_80000_M1 32000_80000_M1 0.020
r 32000_80000_M1 34000_80000_M1 0.020
r 34000_80000_M1 36000_80000_M1 0.020
r 36000_80000_M1 38000_80000_M1 0.020
r 38000_80000_M1 40000_80000_M1 0.020
r 40000_80000_M1 42000_80000_M1 0.020
r 42000_80000_M1 44000_80000_M1 0.020
r 44000_80000_M1 46000_80000_M1 0.020
r 46000_80000_M1 48000_80000_M1 0.020
r 48000_80000_M1 50000_80000_M1 0.020
r 50000_80000_M1 52000_80000_M1 0.020
r 52000_80000_M1 54000_80000_M1 0.020
r 54000_80000_M1 56000_80000_M1 0.020
r 56000_80000_M1 58000_80000_M1 0.020
r 58000_80000_M1 60000_80000_M1 0.020
r 60000_80000_M1 62000_80000_M1 0.020
r 62000_80000_M1 64000_80000_M1 0.020
r 64000_80000_M1 66000_80000_M1 0.020
r 66000_80000_M1 68000_80000_M1 0.020
r 68000_80000_M1 70000_80000_M1 0.020
r 70000_80000_M1 72000_80000_M1 0.020
r 72000_80000_M1 74000_80000_M1 0.020
r 74000_80000_M1 76000_80000_M1 0.020
r 76000_80000_M1 78000_80000_M1 0.020
r 78000_80000_M1 80000_80000_M1 0.020
r 80000_80000_M1 82000_80000_M1 0.020
r 82000_80000_M1 84000_80000_M1 0.020
r 84000_80000_M1 86000_80000_M1 0.020
r 86000_80000_M1 88000_80000_M1 0.020
r 88000_80000_M1 90000_80000_M1 0.020
r 90000_80000_M1 92000_80000_M1 0.020
r 92000_80000_M1 94000_80000_M1 0.020
r 94000_80000_M1 96000_80000_M1 0.020
r 96000_80000_M1 98000_80000_M1 0.020
r 98000_80000_M1 100000_80000_M1 0.020
r 2000_82000_M1 4000_82000_M1 0.020
r 4000_82000_M1 6000_82000_M1 0.020
r 6000_82000_M1 8000_82000_M1 0.020
r 8000_82000_M1 10000_82000_M1 0.020
r 10000_82000_M1 12000_82000_M1 0.020
r 12000_82000_M1 14000_82000_M1 0.020
r 14000_82000_M1 16000_82000_M1 0.020
r 16000_82000_M1 18000_82000_M1 0.020
r 18000_82000_M1 20000_82000_M1 0.020
r 20000_82000_M1 22000_82000_M1 0.020
r 22000_82000_M1 24000_82000_M1 0.020
r 24000_82000_M1 26000_82000_M1 0.020
r 26000_82000_M1 28000_82000_M1 0.020
r 28000_82000_M1 30000_82000_M1 0.020
r 30000_82000_M1 32000_82000_M1 0.020
r 32000_82000_M1 34000_82000_M1 0.020
r 34000_82000_M1 36000_82000_M1 0.020
r 36000_82000_M1 38000_82000_M1 0.020
r 38000_82000_M1 40000_82000_M1 0.020
r 40000_82000_M1 42000_82000_M1 0.020
r 42000_82000_M1 44000_82000_M1 0.020
r 44000_82000_M1 46000_82000_M1 0.020
r 46000_82000_M1 48000_82000_M1 0.020
r 48000_82000_M1 50000_82000_M1 0.020
r 50000_82000_M1 52000_82000_M1 0.020
r 52000_82000_M1 54000_82000_M1 0.020
r 54000_82000_M1 56000_82000_M1 0.020
r 56000_82000_M1 58000_82000_M1 0.020
r 58000_82000_M1 60000_82000_M1 0.020
r 60000_82000_M1 62000_82000_M1 0.020
r 62000_82000_M1 64000_82000_M1 0.020
r 64000_82000_M1 66000_82000_M1 0.020
r 66000_82000_M1 68000_82000_M1 0.020
r 68000_82000_M1 70000_82000_M1 0.020
r 70000_82000_M1 72000_82000_M1 0.020
r 72000_82000_M1 74000_82000_M1 0.020
r 74000_82000_M1 76000_82000_M1 0.020
r 76000_82000_M1 78000_82000_M1 0.020
r 78000_82000_M1 80000_82000_M1 0.020
r 80000_82000_M1 82000_82000_M1 0.020
r 82000_82000_M1 84000_82000_M1 0.020
r 84000_82000_M1 86000_82000_M1 0.020
r 86000_82000_M1 88000_82000_M1 0.020
r 88000_82000_M1 90000_82000_M1 0.020
r 90000_82000_M1 92000_82000_M1 0.020
r 92000_82000_M1 94000_82000_M1 0.020
r 94000_82000_M1 96000_82000_M1 0.020
r 96000_82000_M1 98000_82000_M1 0.020
r 98000_82000_M1 100000_82000_M1 0.020
r 2000_84000_M1 4000_84000_M1 0.020
r 4000_84000_M1 6000_84000_M1 0.020
r 6000_84000_M1 8000_84000_M1 0.020
r 8000_84000_M1 10000_84000_M1 0.020
r 10000_84000_M1 12000_84000_M1 0.020
r 12000_84000_M1 14000_84000_M1 0.020
r 14000_84000_M1 16000_84000_M1 0.020
r 16000_84000_M1 18000_84000_M1 0.020
r 18000_84000_M1 20000_84000_M1 0.020
r 20000_84000_M1 22000_84000_M1 0.020
r 22000_84000_M1 24000_84000_M1 0.020
r 24000_84000_M1 26000_84000_M1 0.020
r 26000_84000_M1 28000_84000_M1 0.020
r 28000_84000_M1 30000_84000_M1 0.020
r 30000_84000_M1 32000_84000_M1 0.020
r 32000_84000_M1 34000_84000_M1 0.020
r 34000_84000_M1 36000_84000_M1 0.020
r 36000_84000_M1 38000_84000_M1 0.020
r 38000_84000_M1 40000_84000_M1 0.020
r 40000_84000_M1 42000_84000_M1 0.020
r 42000_84000_M1 44000_84000_M1 0.020
r 44000_84000_M1 46000_84000_M1 0.020
r 46000_84000_M1 48000_84000_M1 0.020
r 48000_84000_M1 50000_84000_M1 0.020
r 50000_84000_M1 52000_84000_M1 0.020
r 52000_84000_M1 54000_84000_M1 0.020
r 54000_84000_M1 56000_84000_M1 0.020
r 56000_84000_M1 58000_84000_M1 0.020
r 58000_84000_M1 60000_84000_M1 0.020
r 60000_84000_M1 62000_84000_M1 0.020
r 62000_84000_M1 64000_84000_M1 0.020
r 64000_84000_M1 66000_84000_M1 0.020
r 66000_84000_M1 68000_84000_M1 0.020
r 68000_84000_M1 70000_84000_M1 0.020
r 70000_84000_M1 72000_84000_M1 0.020
r 72000_84000_M1 74000_84000_M1 0.020
r 74000_84000_M1 76000_84000_M1 0.020
r 76000_84000_M1 78000_84000_M1 0.020
r 78000_84000_M1 80000_84000_M1 0.020
r 80000_84000_M1 82000_84000_M1 0.020
r 82000_84000_M1 84000_84000_M1 0.020
r 84000_84000_M1 86000_84000_M1 0.020
r 86000_84000_M1 88000_84000_M1 0.020
r 88000_84000_M1 90000_84000_M1 0.020
r 90000_84000_M1 92000_84000_M1 0.020
r 92000_84000_M1 94000_84000_M1 0.020
r 94000_84000_M1 96000_84000_M1 0.020
r 96000_84000_M1 98000_84000_M1 0.020
r 98000_84000_M1 100000_84000_M1 0.020
r 2000_86000_M1 4000_86000_M1 0.020
r 4000_86000_M1 6000_86000_M1 0.020
r 6000_86000_M1 8000_86000_M1 0.020
r 8000_86000_M1 10000_86000_M1 0.020
r 10000_86000_M1 12000_86000_M1 0.020
r 12000_86000_M1 14000_86000_M1 0.020
r 14000_86000_M1 16000_86000_M1 0.020
r 16000_86000_M1 18000_86000_M1 0.020
r 18000_86000_M1 20000_86000_M1 0.020
r 20000_86000_M1 22000_86000_M1 0.020
r 22000_86000_M1 24000_86000_M1 0.020
r 24000_86000_M1 26000_86000_M1 0.020
r 26000_86000_M1 28000_86000_M1 0.020
r 28000_86000_M1 30000_86000_M1 0.020
r 30000_86000_M1 32000_86000_M1 0.020
r 32000_86000_M1 34000_86000_M1 0.020
r 34000_86000_M1 36000_86000_M1 0.020
r 36000_86000_M1 38000_86000_M1 0.020
r 38000_86000_M1 40000_86000_M1 0.020
r 40000_86000_M1 42000_86000_M1 0.020
r 42000_86000_M1 44000_86000_M1 0.020
r 44000_86000_M1 46000_86000_M1 0.020
r 46000_86000_M1 48000_86000_M1 0.020
r 48000_86000_M1 50000_86000_M1 0.020
r 50000_86000_M1 52000_86000_M1 0.020
r 52000_86000_M1 54000_86000_M1 0.020
r 54000_86000_M1 56000_86000_M1 0.020
r 56000_86000_M1 58000_86000_M1 0.020
r 58000_86000_M1 60000_86000_M1 0.020
r 60000_86000_M1 62000_86000_M1 0.020
r 62000_86000_M1 64000_86000_M1 0.020
r 64000_86000_M1 66000_86000_M1 0.020
r 66000_86000_M1 68000_86000_M1 0.020
r 68000_86000_M1 70000_86000_M1 0.020
r 70000_86000_M1 72000_86000_M1 0.020
r 72000_86000_M1 74000_86000_M1 0.020
r 74000_86000_M1 76000_86000_M1 0.020
r 76000_86000_M1 78000_86000_M1 0.020
r 78000_86000_M1 80000_86000_M1 0.020
r 80000_86000_M1 82000_86000_M1 0.020
r 82000_86000_M1 84000_86000_M1 0.020
r 84000_86000_M1 86000_86000_M1 0.020
r 86000_86000_M1 88000_86000_M1 0.020
r 88000_86000_M1 90000_86000_M1 0.020
r 90000_86000_M1 92000_86000_M1 0.020
r 92000_86000_M1 94000_86000_M1 0.020
r 94000_86000_M1 96000_86000_M1 0.020
r 96000_86000_M1 98000_86000_M1 0.020
r 98000_86000_M1 100000_86000_M1 0.020
r 2000_88000_M1 4000_88000_M1 0.020
r 4000_88000_M1 6000_88000_M1 0.020
r 6000_88000_M1 8000_88000_M1 0.020
r 8000_88000_M1 10000_88000_M1 0.020
r 10000_88000_M1 12000_88000_M1 0.020
r 12000_88000_M1 14000_88000_M1 0.020
r 14000_88000_M1 16000_88000_M1 0.020
r 16000_88000_M1 18000_88000_M1 0.020
r 18000_88000_M1 20000_88000_M1 0.020
r 20000_88000_M1 22000_88000_M1 0.020
r 22000_88000_M1 24000_88000_M1 0.020
r 24000_88000_M1 26000_88000_M1 0.020
r 26000_88000_M1 28000_88000_M1 0.020
r 28000_88000_M1 30000_88000_M1 0.020
r 30000_88000_M1 32000_88000_M1 0.020
r 32000_88000_M1 34000_88000_M1 0.020
r 34000_88000_M1 36000_88000_M1 0.020
r 36000_88000_M1 38000_88000_M1 0.020
r 38000_88000_M1 40000_88000_M1 0.020
r 40000_88000_M1 42000_88000_M1 0.020
r 42000_88000_M1 44000_88000_M1 0.020
r 44000_88000_M1 46000_88000_M1 0.020
r 46000_88000_M1 48000_88000_M1 0.020
r 48000_88000_M1 50000_88000_M1 0.020
r 50000_88000_M1 52000_88000_M1 0.020
r 52000_88000_M1 54000_88000_M1 0.020
r 54000_88000_M1 56000_88000_M1 0.020
r 56000_88000_M1 58000_88000_M1 0.020
r 58000_88000_M1 60000_88000_M1 0.020
r 60000_88000_M1 62000_88000_M1 0.020
r 62000_88000_M1 64000_88000_M1 0.020
r 64000_88000_M1 66000_88000_M1 0.020
r 66000_88000_M1 68000_88000_M1 0.020
r 68000_88000_M1 70000_88000_M1 0.020
r 70000_88000_M1 72000_88000_M1 0.020
r 72000_88000_M1 74000_88000_M1 0.020
r 74000_88000_M1 76000_88000_M1 0.020
r 76000_88000_M1 78000_88000_M1 0.020
r 78000_88000_M1 80000_88000_M1 0.020
r 80000_88000_M1 82000_88000_M1 0.020
r 82000_88000_M1 84000_88000_M1 0.020
r 84000_88000_M1 86000_88000_M1 0.020
r 86000_88000_M1 88000_88000_M1 0.020
r 88000_88000_M1 90000_88000_M1 0.020
r 90000_88000_M1 92000_88000_M1 0.020
r 92000_88000_M1 94000_88000_M1 0.020
r 94000_88000_M1 96000_88000_M1 0.020
r 96000_88000_M1 98000_88000_M1 0.020
r 98000_88000_M1 100000_88000_M1 0.020
r 2000_90000_M1 4000_90000_M1 0.020
r 4000_90000_M1 6000_90000_M1 0.020
r 6000_90000_M1 8000_90000_M1 0.020
r 8000_90000_M1 10000_90000_M1 0.020
r 10000_90000_M1 12000_90000_M1 0.020
r 12000_90000_M1 14000_90000_M1 0.020
r 14000_90000_M1 16000_90000_M1 0.020
r 16000_90000_M1 18000_90000_M1 0.020
r 18000_90000_M1 20000_90000_M1 0.020
r 20000_90000_M1 22000_90000_M1 0.020
r 22000_90000_M1 24000_90000_M1 0.020
r 24000_90000_M1 26000_90000_M1 0.020
r 26000_90000_M1 28000_90000_M1 0.020
r 28000_90000_M1 30000_90000_M1 0.020
r 30000_90000_M1 32000_90000_M1 0.020
r 32000_90000_M1 34000_90000_M1 0.020
r 34000_90000_M1 36000_90000_M1 0.020
r 36000_90000_M1 38000_90000_M1 0.020
r 38000_90000_M1 40000_90000_M1 0.020
r 40000_90000_M1 42000_90000_M1 0.020
r 42000_90000_M1 44000_90000_M1 0.020
r 44000_90000_M1 46000_90000_M1 0.020
r 46000_90000_M1 48000_90000_M1 0.020
r 48000_90000_M1 50000_90000_M1 0.020
r 50000_90000_M1 52000_90000_M1 0.020
r 52000_90000_M1 54000_90000_M1 0.020
r 54000_90000_M1 56000_90000_M1 0.020
r 56000_90000_M1 58000_90000_M1 0.020
r 58000_90000_M1 60000_90000_M1 0.020
r 60000_90000_M1 62000_90000_M1 0.020
r 62000_90000_M1 64000_90000_M1 0.020
r 64000_90000_M1 66000_90000_M1 0.020
r 66000_90000_M1 68000_90000_M1 0.020
r 68000_90000_M1 70000_90000_M1 0.020
r 70000_90000_M1 72000_90000_M1 0.020
r 72000_90000_M1 74000_90000_M1 0.020
r 74000_90000_M1 76000_90000_M1 0.020
r 76000_90000_M1 78000_90000_M1 0.020
r 78000_90000_M1 80000_90000_M1 0.020
r 80000_90000_M1 82000_90000_M1 0.020
r 82000_90000_M1 84000_90000_M1 0.020
r 84000_90000_M1 86000_90000_M1 0.020
r 86000_90000_M1 88000_90000_M1 0.020
r 88000_90000_M1 90000_90000_M1 0.020
r 90000_90000_M1 92000_90000_M1 0.020
r 92000_90000_M1 94000_90000_M1 0.020
r 94000_90000_M1 96000_90000_M1 0.020
r 96000_90000_M1 98000_90000_M1 0.020
r 98000_90000_M1 100000_90000_M1 0.020
r 2000_92000_M1 4000_92000_M1 0.020
r 4000_92000_M1 6000_92000_M1 0.020
r 6000_92000_M1 8000_92000_M1 0.020
r 8000_92000_M1 10000_92000_M1 0.020
r 10000_92000_M1 12000_92000_M1 0.020
r 12000_92000_M1 14000_92000_M1 0.020
r 14000_92000_M1 16000_92000_M1 0.020
r 16000_92000_M1 18000_92000_M1 0.020
r 18000_92000_M1 20000_92000_M1 0.020
r 20000_92000_M1 22000_92000_M1 0.020
r 22000_92000_M1 24000_92000_M1 0.020
r 24000_92000_M1 26000_92000_M1 0.020
r 26000_92000_M1 28000_92000_M1 0.020
r 28000_92000_M1 30000_92000_M1 0.020
r 30000_92000_M1 32000_92000_M1 0.020
r 32000_92000_M1 34000_92000_M1 0.020
r 34000_92000_M1 36000_92000_M1 0.020
r 36000_92000_M1 38000_92000_M1 0.020
r 38000_92000_M1 40000_92000_M1 0.020
r 40000_92000_M1 42000_92000_M1 0.020
r 42000_92000_M1 44000_92000_M1 0.020
r 44000_92000_M1 46000_92000_M1 0.020
r 46000_92000_M1 48000_92000_M1 0.020
r 48000_92000_M1 50000_92000_M1 0.020
r 50000_92000_M1 52000_92000_M1 0.020
r 52000_92000_M1 54000_92000_M1 0.020
r 54000_92000_M1 56000_92000_M1 0.020
r 56000_92000_M1 58000_92000_M1 0.020
r 58000_92000_M1 60000_92000_M1 0.020
r 60000_92000_M1 62000_92000_M1 0.020
r 62000_92000_M1 64000_92000_M1 0.020
r 64000_92000_M1 66000_92000_M1 0.020
r 66000_92000_M1 68000_92000_M1 0.020
r 68000_92000_M1 70000_92000_M1 0.020
r 70000_92000_M1 72000_92000_M1 0.020
r 72000_92000_M1 74000_92000_M1 0.020
r 74000_92000_M1 76000_92000_M1 0.020
r 76000_92000_M1 78000_92000_M1 0.020
r 78000_92000_M1 80000_92000_M1 0.020
r 80000_92000_M1 82000_92000_M1 0.020
r 82000_92000_M1 84000_92000_M1 0.020
r 84000_92000_M1 86000_92000_M1 0.020
r 86000_92000_M1 88000_92000_M1 0.020
r 88000_92000_M1 90000_92000_M1 0.020
r 90000_92000_M1 92000_92000_M1 0.020
r 92000_92000_M1 94000_92000_M1 0.020
r 94000_92000_M1 96000_92000_M1 0.020
r 96000_92000_M1 98000_92000_M1 0.020
r 98000_92000_M1 100000_92000_M1 0.020
r 2000_94000_M1 4000_94000_M1 0.020
r 4000_94000_M1 6000_94000_M1 0.020
r 6000_94000_M1 8000_94000_M1 0.020
r 8000_94000_M1 10000_94000_M1 0.020
r 10000_94000_M1 12000_94000_M1 0.020
r 12000_94000_M1 14000_94000_M1 0.020
r 14000_94000_M1 16000_94000_M1 0.020
r 16000_94000_M1 18000_94000_M1 0.020
r 18000_94000_M1 20000_94000_M1 0.020
r 20000_94000_M1 22000_94000_M1 0.020
r 22000_94000_M1 24000_94000_M1 0.020
r 24000_94000_M1 26000_94000_M1 0.020
r 26000_94000_M1 28000_94000_M1 0.020
r 28000_94000_M1 30000_94000_M1 0.020
r 30000_94000_M1 32000_94000_M1 0.020
r 32000_94000_M1 34000_94000_M1 0.020
r 34000_94000_M1 36000_94000_M1 0.020
r 36000_94000_M1 38000_94000_M1 0.020
r 38000_94000_M1 40000_94000_M1 0.020
r 40000_94000_M1 42000_94000_M1 0.020
r 42000_94000_M1 44000_94000_M1 0.020
r 44000_94000_M1 46000_94000_M1 0.020
r 46000_94000_M1 48000_94000_M1 0.020
r 48000_94000_M1 50000_94000_M1 0.020
r 50000_94000_M1 52000_94000_M1 0.020
r 52000_94000_M1 54000_94000_M1 0.020
r 54000_94000_M1 56000_94000_M1 0.020
r 56000_94000_M1 58000_94000_M1 0.020
r 58000_94000_M1 60000_94000_M1 0.020
r 60000_94000_M1 62000_94000_M1 0.020
r 62000_94000_M1 64000_94000_M1 0.020
r 64000_94000_M1 66000_94000_M1 0.020
r 66000_94000_M1 68000_94000_M1 0.020
r 68000_94000_M1 70000_94000_M1 0.020
r 70000_94000_M1 72000_94000_M1 0.020
r 72000_94000_M1 74000_94000_M1 0.020
r 74000_94000_M1 76000_94000_M1 0.020
r 76000_94000_M1 78000_94000_M1 0.020
r 78000_94000_M1 80000_94000_M1 0.020
r 80000_94000_M1 82000_94000_M1 0.020
r 82000_94000_M1 84000_94000_M1 0.020
r 84000_94000_M1 86000_94000_M1 0.020
r 86000_94000_M1 88000_94000_M1 0.020
r 88000_94000_M1 90000_94000_M1 0.020
r 90000_94000_M1 92000_94000_M1 0.020
r 92000_94000_M1 94000_94000_M1 0.020
r 94000_94000_M1 96000_94000_M1 0.020
r 96000_94000_M1 98000_94000_M1 0.020
r 98000_94000_M1 100000_94000_M1 0.020
r 2000_96000_M1 4000_96000_M1 0.020
r 4000_96000_M1 6000_96000_M1 0.020
r 6000_96000_M1 8000_96000_M1 0.020
r 8000_96000_M1 10000_96000_M1 0.020
r 10000_96000_M1 12000_96000_M1 0.020
r 12000_96000_M1 14000_96000_M1 0.020
r 14000_96000_M1 16000_96000_M1 0.020
r 16000_96000_M1 18000_96000_M1 0.020
r 18000_96000_M1 20000_96000_M1 0.020
r 20000_96000_M1 22000_96000_M1 0.020
r 22000_96000_M1 24000_96000_M1 0.020
r 24000_96000_M1 26000_96000_M1 0.020
r 26000_96000_M1 28000_96000_M1 0.020
r 28000_96000_M1 30000_96000_M1 0.020
r 30000_96000_M1 32000_96000_M1 0.020
r 32000_96000_M1 34000_96000_M1 0.020
r 34000_96000_M1 36000_96000_M1 0.020
r 36000_96000_M1 38000_96000_M1 0.020
r 38000_96000_M1 40000_96000_M1 0.020
r 40000_96000_M1 42000_96000_M1 0.020
r 42000_96000_M1 44000_96000_M1 0.020
r 44000_96000_M1 46000_96000_M1 0.020
r 46000_96000_M1 48000_96000_M1 0.020
r 48000_96000_M1 50000_96000_M1 0.020
r 50000_96000_M1 52000_96000_M1 0.020
r 52000_96000_M1 54000_96000_M1 0.020
r 54000_96000_M1 56000_96000_M1 0.020
r 56000_96000_M1 58000_96000_M1 0.020
r 58000_96000_M1 60000_96000_M1 0.020
r 60000_96000_M1 62000_96000_M1 0.020
r 62000_96000_M1 64000_96000_M1 0.020
r 64000_96000_M1 66000_96000_M1 0.020
r 66000_96000_M1 68000_96000_M1 0.020
r 68000_96000_M1 70000_96000_M1 0.020
r 70000_96000_M1 72000_96000_M1 0.020
r 72000_96000_M1 74000_96000_M1 0.020
r 74000_96000_M1 76000_96000_M1 0.020
r 76000_96000_M1 78000_96000_M1 0.020
r 78000_96000_M1 80000_96000_M1 0.020
r 80000_96000_M1 82000_96000_M1 0.020
r 82000_96000_M1 84000_96000_M1 0.020
r 84000_96000_M1 86000_96000_M1 0.020
r 86000_96000_M1 88000_96000_M1 0.020
r 88000_96000_M1 90000_96000_M1 0.020
r 90000_96000_M1 92000_96000_M1 0.020
r 92000_96000_M1 94000_96000_M1 0.020
r 94000_96000_M1 96000_96000_M1 0.020
r 96000_96000_M1 98000_96000_M1 0.020
r 98000_96000_M1 100000_96000_M1 0.020
r 2000_98000_M1 4000_98000_M1 0.020
r 4000_98000_M1 6000_98000_M1 0.020
r 6000_98000_M1 8000_98000_M1 0.020
r 8000_98000_M1 10000_98000_M1 0.020
r 10000_98000_M1 12000_98000_M1 0.020
r 12000_98000_M1 14000_98000_M1 0.020
r 14000_98000_M1 16000_98000_M1 0.020
r 16000_98000_M1 18000_98000_M1 0.020
r 18000_98000_M1 20000_98000_M1 0.020
r 20000_98000_M1 22000_98000_M1 0.020
r 22000_98000_M1 24000_98000_M1 0.020
r 24000_98000_M1 26000_98000_M1 0.020
r 26000_98000_M1 28000_98000_M1 0.020
r 28000_98000_M1 30000_98000_M1 0.020
r 30000_98000_M1 32000_98000_M1 0.020
r 32000_98000_M1 34000_98000_M1 0.020
r 34000_98000_M1 36000_98000_M1 0.020
r 36000_98000_M1 38000_98000_M1 0.020
r 38000_98000_M1 40000_98000_M1 0.020
r 40000_98000_M1 42000_98000_M1 0.020
r 42000_98000_M1 44000_98000_M1 0.020
r 44000_98000_M1 46000_98000_M1 0.020
r 46000_98000_M1 48000_98000_M1 0.020
r 48000_98000_M1 50000_98000_M1 0.020
r 50000_98000_M1 52000_98000_M1 0.020
r 52000_98000_M1 54000_98000_M1 0.020
r 54000_98000_M1 56000_98000_M1 0.020
r 56000_98000_M1 58000_98000_M1 0.020
r 58000_98000_M1 60000_98000_M1 0.020
r 60000_98000_M1 62000_98000_M1 0.020
r 62000_98000_M1 64000_98000_M1 0.020
r 64000_98000_M1 66000_98000_M1 0.020
r 66000_98000_M1 68000_98000_M1 0.020
r 68000_98000_M1 70000_98000_M1 0.020
r 70000_98000_M1 72000_98000_M1 0.020
r 72000_98000_M1 74000_98000_M1 0.020
r 74000_98000_M1 76000_98000_M1 0.020
r 76000_98000_M1 78000_98000_M1 0.020
r 78000_98000_M1 80000_98000_M1 0.020
r 80000_98000_M1 82000_98000_M1 0.020
r 82000_98000_M1 84000_98000_M1 0.020
r 84000_98000_M1 86000_98000_M1 0.020
r 86000_98000_M1 88000_98000_M1 0.020
r 88000_98000_M1 90000_98000_M1 0.020
r 90000_98000_M1 92000_98000_M1 0.020
r 92000_98000_M1 94000_98000_M1 0.020
r 94000_98000_M1 96000_98000_M1 0.020
r 96000_98000_M1 98000_98000_M1 0.020
r 98000_98000_M1 100000_98000_M1 0.020
r 2000_100000_M1 4000_100000_M1 0.020
r 4000_100000_M1 6000_100000_M1 0.020
r 6000_100000_M1 8000_100000_M1 0.020
r 8000_100000_M1 10000_100000_M1 0.020
r 10000_100000_M1 12000_100000_M1 0.020
r 12000_100000_M1 14000_100000_M1 0.020
r 14000_100000_M1 16000_100000_M1 0.020
r 16000_100000_M1 18000_100000_M1 0.020
r 18000_100000_M1 20000_100000_M1 0.020
r 20000_100000_M1 22000_100000_M1 0.020
r 22000_100000_M1 24000_100000_M1 0.020
r 24000_100000_M1 26000_100000_M1 0.020
r 26000_100000_M1 28000_100000_M1 0.020
r 28000_100000_M1 30000_100000_M1 0.020
r 30000_100000_M1 32000_100000_M1 0.020
r 32000_100000_M1 34000_100000_M1 0.020
r 34000_100000_M1 36000_100000_M1 0.020
r 36000_100000_M1 38000_100000_M1 0.020
r 38000_100000_M1 40000_100000_M1 0.020
r 40000_100000_M1 42000_100000_M1 0.020
r 42000_100000_M1 44000_100000_M1 0.020
r 44000_100000_M1 46000_100000_M1 0.020
r 46000_100000_M1 48000_100000_M1 0.020
r 48000_100000_M1 50000_100000_M1 0.020
r 50000_100000_M1 52000_100000_M1 0.020
r 52000_100000_M1 54000_100000_M1 0.020
r 54000_100000_M1 56000_100000_M1 0.020
r 56000_100000_M1 58000_100000_M1 0.020
r 58000_100000_M1 60000_100000_M1 0.020
r 60000_100000_M1 62000_100000_M1 0.020
r 62000_100000_M1 64000_100000_M1 0.020
r 64000_100000_M1 66000_100000_M1 0.020
r 66000_100000_M1 68000_100000_M1 0.020
r 68000_100000_M1 70000_100000_M1 0.020
r 70000_100000_M1 72000_100000_M1 0.020
r 72000_100000_M1 74000_100000_M1 0.020
r 74000_100000_M1 76000_100000_M1 0.020
r 76000_100000_M1 78000_100000_M1 0.020
r 78000_100000_M1 80000_100000_M1 0.020
r 80000_100000_M1 82000_100000_M1 0.020
r 82000_100000_M1 84000_100000_M1 0.020
r 84000_100000_M1 86000_100000_M1 0.020
r 86000_100000_M1 88000_100000_M1 0.020
r 88000_100000_M1 90000_100000_M1 0.020
r 90000_100000_M1 92000_100000_M1 0.020
r 92000_100000_M1 94000_100000_M1 0.020
r 94000_100000_M1 96000_100000_M1 0.020
r 96000_100000_M1 98000_100000_M1 0.020
r 98000_100000_M1 100000_100000_M1 0.020

* M1 Vertical resistors
r 2000_2000_M1 2000_4000_M1 0.025
r 2000_4000_M1 2000_6000_M1 0.025
r 2000_6000_M1 2000_8000_M1 0.025
r 2000_8000_M1 2000_10000_M1 0.025
r 2000_10000_M1 2000_12000_M1 0.025
r 2000_12000_M1 2000_14000_M1 0.025
r 2000_14000_M1 2000_16000_M1 0.025
r 2000_16000_M1 2000_18000_M1 0.025
r 2000_18000_M1 2000_20000_M1 0.025
r 2000_20000_M1 2000_22000_M1 0.025
r 2000_22000_M1 2000_24000_M1 0.025
r 2000_24000_M1 2000_26000_M1 0.025
r 2000_26000_M1 2000_28000_M1 0.025
r 2000_28000_M1 2000_30000_M1 0.025
r 2000_30000_M1 2000_32000_M1 0.025
r 2000_32000_M1 2000_34000_M1 0.025
r 2000_34000_M1 2000_36000_M1 0.025
r 2000_36000_M1 2000_38000_M1 0.025
r 2000_38000_M1 2000_40000_M1 0.025
r 2000_40000_M1 2000_42000_M1 0.025
r 2000_42000_M1 2000_44000_M1 0.025
r 2000_44000_M1 2000_46000_M1 0.025
r 2000_46000_M1 2000_48000_M1 0.025
r 2000_48000_M1 2000_50000_M1 0.025
r 2000_50000_M1 2000_52000_M1 0.025
r 2000_52000_M1 2000_54000_M1 0.025
r 2000_54000_M1 2000_56000_M1 0.025
r 2000_56000_M1 2000_58000_M1 0.025
r 2000_58000_M1 2000_60000_M1 0.025
r 2000_60000_M1 2000_62000_M1 0.025
r 2000_62000_M1 2000_64000_M1 0.025
r 2000_64000_M1 2000_66000_M1 0.025
r 2000_66000_M1 2000_68000_M1 0.025
r 2000_68000_M1 2000_70000_M1 0.025
r 2000_70000_M1 2000_72000_M1 0.025
r 2000_72000_M1 2000_74000_M1 0.025
r 2000_74000_M1 2000_76000_M1 0.025
r 2000_76000_M1 2000_78000_M1 0.025
r 2000_78000_M1 2000_80000_M1 0.025
r 2000_80000_M1 2000_82000_M1 0.025
r 2000_82000_M1 2000_84000_M1 0.025
r 2000_84000_M1 2000_86000_M1 0.025
r 2000_86000_M1 2000_88000_M1 0.025
r 2000_88000_M1 2000_90000_M1 0.025
r 2000_90000_M1 2000_92000_M1 0.025
r 2000_92000_M1 2000_94000_M1 0.025
r 2000_94000_M1 2000_96000_M1 0.025
r 2000_96000_M1 2000_98000_M1 0.025
r 2000_98000_M1 2000_100000_M1 0.025
r 4000_2000_M1 4000_4000_M1 0.025
r 4000_4000_M1 4000_6000_M1 0.025
r 4000_6000_M1 4000_8000_M1 0.025
r 4000_8000_M1 4000_10000_M1 0.025
r 4000_10000_M1 4000_12000_M1 0.025
r 4000_12000_M1 4000_14000_M1 0.025
r 4000_14000_M1 4000_16000_M1 0.025
r 4000_16000_M1 4000_18000_M1 0.025
r 4000_18000_M1 4000_20000_M1 0.025
r 4000_20000_M1 4000_22000_M1 0.025
r 4000_22000_M1 4000_24000_M1 0.025
r 4000_24000_M1 4000_26000_M1 0.025
r 4000_26000_M1 4000_28000_M1 0.025
r 4000_28000_M1 4000_30000_M1 0.025
r 4000_30000_M1 4000_32000_M1 0.025
r 4000_32000_M1 4000_34000_M1 0.025
r 4000_34000_M1 4000_36000_M1 0.025
r 4000_36000_M1 4000_38000_M1 0.025
r 4000_38000_M1 4000_40000_M1 0.025
r 4000_40000_M1 4000_42000_M1 0.025
r 4000_42000_M1 4000_44000_M1 0.025
r 4000_44000_M1 4000_46000_M1 0.025
r 4000_46000_M1 4000_48000_M1 0.025
r 4000_48000_M1 4000_50000_M1 0.025
r 4000_50000_M1 4000_52000_M1 0.025
r 4000_52000_M1 4000_54000_M1 0.025
r 4000_54000_M1 4000_56000_M1 0.025
r 4000_56000_M1 4000_58000_M1 0.025
r 4000_58000_M1 4000_60000_M1 0.025
r 4000_60000_M1 4000_62000_M1 0.025
r 4000_62000_M1 4000_64000_M1 0.025
r 4000_64000_M1 4000_66000_M1 0.025
r 4000_66000_M1 4000_68000_M1 0.025
r 4000_68000_M1 4000_70000_M1 0.025
r 4000_70000_M1 4000_72000_M1 0.025
r 4000_72000_M1 4000_74000_M1 0.025
r 4000_74000_M1 4000_76000_M1 0.025
r 4000_76000_M1 4000_78000_M1 0.025
r 4000_78000_M1 4000_80000_M1 0.025
r 4000_80000_M1 4000_82000_M1 0.025
r 4000_82000_M1 4000_84000_M1 0.025
r 4000_84000_M1 4000_86000_M1 0.025
r 4000_86000_M1 4000_88000_M1 0.025
r 4000_88000_M1 4000_90000_M1 0.025
r 4000_90000_M1 4000_92000_M1 0.025
r 4000_92000_M1 4000_94000_M1 0.025
r 4000_94000_M1 4000_96000_M1 0.025
r 4000_96000_M1 4000_98000_M1 0.025
r 4000_98000_M1 4000_100000_M1 0.025
r 6000_2000_M1 6000_4000_M1 0.025
r 6000_4000_M1 6000_6000_M1 0.025
r 6000_6000_M1 6000_8000_M1 0.025
r 6000_8000_M1 6000_10000_M1 0.025
r 6000_10000_M1 6000_12000_M1 0.025
r 6000_12000_M1 6000_14000_M1 0.025
r 6000_14000_M1 6000_16000_M1 0.025
r 6000_16000_M1 6000_18000_M1 0.025
r 6000_18000_M1 6000_20000_M1 0.025
r 6000_20000_M1 6000_22000_M1 0.025
r 6000_22000_M1 6000_24000_M1 0.025
r 6000_24000_M1 6000_26000_M1 0.025
r 6000_26000_M1 6000_28000_M1 0.025
r 6000_28000_M1 6000_30000_M1 0.025
r 6000_30000_M1 6000_32000_M1 0.025
r 6000_32000_M1 6000_34000_M1 0.025
r 6000_34000_M1 6000_36000_M1 0.025
r 6000_36000_M1 6000_38000_M1 0.025
r 6000_38000_M1 6000_40000_M1 0.025
r 6000_40000_M1 6000_42000_M1 0.025
r 6000_42000_M1 6000_44000_M1 0.025
r 6000_44000_M1 6000_46000_M1 0.025
r 6000_46000_M1 6000_48000_M1 0.025
r 6000_48000_M1 6000_50000_M1 0.025
r 6000_50000_M1 6000_52000_M1 0.025
r 6000_52000_M1 6000_54000_M1 0.025
r 6000_54000_M1 6000_56000_M1 0.025
r 6000_56000_M1 6000_58000_M1 0.025
r 6000_58000_M1 6000_60000_M1 0.025
r 6000_60000_M1 6000_62000_M1 0.025
r 6000_62000_M1 6000_64000_M1 0.025
r 6000_64000_M1 6000_66000_M1 0.025
r 6000_66000_M1 6000_68000_M1 0.025
r 6000_68000_M1 6000_70000_M1 0.025
r 6000_70000_M1 6000_72000_M1 0.025
r 6000_72000_M1 6000_74000_M1 0.025
r 6000_74000_M1 6000_76000_M1 0.025
r 6000_76000_M1 6000_78000_M1 0.025
r 6000_78000_M1 6000_80000_M1 0.025
r 6000_80000_M1 6000_82000_M1 0.025
r 6000_82000_M1 6000_84000_M1 0.025
r 6000_84000_M1 6000_86000_M1 0.025
r 6000_86000_M1 6000_88000_M1 0.025
r 6000_88000_M1 6000_90000_M1 0.025
r 6000_90000_M1 6000_92000_M1 0.025
r 6000_92000_M1 6000_94000_M1 0.025
r 6000_94000_M1 6000_96000_M1 0.025
r 6000_96000_M1 6000_98000_M1 0.025
r 6000_98000_M1 6000_100000_M1 0.025
r 8000_2000_M1 8000_4000_M1 0.025
r 8000_4000_M1 8000_6000_M1 0.025
r 8000_6000_M1 8000_8000_M1 0.025
r 8000_8000_M1 8000_10000_M1 0.025
r 8000_10000_M1 8000_12000_M1 0.025
r 8000_12000_M1 8000_14000_M1 0.025
r 8000_14000_M1 8000_16000_M1 0.025
r 8000_16000_M1 8000_18000_M1 0.025
r 8000_18000_M1 8000_20000_M1 0.025
r 8000_20000_M1 8000_22000_M1 0.025
r 8000_22000_M1 8000_24000_M1 0.025
r 8000_24000_M1 8000_26000_M1 0.025
r 8000_26000_M1 8000_28000_M1 0.025
r 8000_28000_M1 8000_30000_M1 0.025
r 8000_30000_M1 8000_32000_M1 0.025
r 8000_32000_M1 8000_34000_M1 0.025
r 8000_34000_M1 8000_36000_M1 0.025
r 8000_36000_M1 8000_38000_M1 0.025
r 8000_38000_M1 8000_40000_M1 0.025
r 8000_40000_M1 8000_42000_M1 0.025
r 8000_42000_M1 8000_44000_M1 0.025
r 8000_44000_M1 8000_46000_M1 0.025
r 8000_46000_M1 8000_48000_M1 0.025
r 8000_48000_M1 8000_50000_M1 0.025
r 8000_50000_M1 8000_52000_M1 0.025
r 8000_52000_M1 8000_54000_M1 0.025
r 8000_54000_M1 8000_56000_M1 0.025
r 8000_56000_M1 8000_58000_M1 0.025
r 8000_58000_M1 8000_60000_M1 0.025
r 8000_60000_M1 8000_62000_M1 0.025
r 8000_62000_M1 8000_64000_M1 0.025
r 8000_64000_M1 8000_66000_M1 0.025
r 8000_66000_M1 8000_68000_M1 0.025
r 8000_68000_M1 8000_70000_M1 0.025
r 8000_70000_M1 8000_72000_M1 0.025
r 8000_72000_M1 8000_74000_M1 0.025
r 8000_74000_M1 8000_76000_M1 0.025
r 8000_76000_M1 8000_78000_M1 0.025
r 8000_78000_M1 8000_80000_M1 0.025
r 8000_80000_M1 8000_82000_M1 0.025
r 8000_82000_M1 8000_84000_M1 0.025
r 8000_84000_M1 8000_86000_M1 0.025
r 8000_86000_M1 8000_88000_M1 0.025
r 8000_88000_M1 8000_90000_M1 0.025
r 8000_90000_M1 8000_92000_M1 0.025
r 8000_92000_M1 8000_94000_M1 0.025
r 8000_94000_M1 8000_96000_M1 0.025
r 8000_96000_M1 8000_98000_M1 0.025
r 8000_98000_M1 8000_100000_M1 0.025
r 10000_2000_M1 10000_4000_M1 0.025
r 10000_4000_M1 10000_6000_M1 0.025
r 10000_6000_M1 10000_8000_M1 0.025
r 10000_8000_M1 10000_10000_M1 0.025
r 10000_10000_M1 10000_12000_M1 0.025
r 10000_12000_M1 10000_14000_M1 0.025
r 10000_14000_M1 10000_16000_M1 0.025
r 10000_16000_M1 10000_18000_M1 0.025
r 10000_18000_M1 10000_20000_M1 0.025
r 10000_20000_M1 10000_22000_M1 0.025
r 10000_22000_M1 10000_24000_M1 0.025
r 10000_24000_M1 10000_26000_M1 0.025
r 10000_26000_M1 10000_28000_M1 0.025
r 10000_28000_M1 10000_30000_M1 0.025
r 10000_30000_M1 10000_32000_M1 0.025
r 10000_32000_M1 10000_34000_M1 0.025
r 10000_34000_M1 10000_36000_M1 0.025
r 10000_36000_M1 10000_38000_M1 0.025
r 10000_38000_M1 10000_40000_M1 0.025
r 10000_40000_M1 10000_42000_M1 0.025
r 10000_42000_M1 10000_44000_M1 0.025
r 10000_44000_M1 10000_46000_M1 0.025
r 10000_46000_M1 10000_48000_M1 0.025
r 10000_48000_M1 10000_50000_M1 0.025
r 10000_50000_M1 10000_52000_M1 0.025
r 10000_52000_M1 10000_54000_M1 0.025
r 10000_54000_M1 10000_56000_M1 0.025
r 10000_56000_M1 10000_58000_M1 0.025
r 10000_58000_M1 10000_60000_M1 0.025
r 10000_60000_M1 10000_62000_M1 0.025
r 10000_62000_M1 10000_64000_M1 0.025
r 10000_64000_M1 10000_66000_M1 0.025
r 10000_66000_M1 10000_68000_M1 0.025
r 10000_68000_M1 10000_70000_M1 0.025
r 10000_70000_M1 10000_72000_M1 0.025
r 10000_72000_M1 10000_74000_M1 0.025
r 10000_74000_M1 10000_76000_M1 0.025
r 10000_76000_M1 10000_78000_M1 0.025
r 10000_78000_M1 10000_80000_M1 0.025
r 10000_80000_M1 10000_82000_M1 0.025
r 10000_82000_M1 10000_84000_M1 0.025
r 10000_84000_M1 10000_86000_M1 0.025
r 10000_86000_M1 10000_88000_M1 0.025
r 10000_88000_M1 10000_90000_M1 0.025
r 10000_90000_M1 10000_92000_M1 0.025
r 10000_92000_M1 10000_94000_M1 0.025
r 10000_94000_M1 10000_96000_M1 0.025
r 10000_96000_M1 10000_98000_M1 0.025
r 10000_98000_M1 10000_100000_M1 0.025
r 12000_2000_M1 12000_4000_M1 0.025
r 12000_4000_M1 12000_6000_M1 0.025
r 12000_6000_M1 12000_8000_M1 0.025
r 12000_8000_M1 12000_10000_M1 0.025
r 12000_10000_M1 12000_12000_M1 0.025
r 12000_12000_M1 12000_14000_M1 0.025
r 12000_14000_M1 12000_16000_M1 0.025
r 12000_16000_M1 12000_18000_M1 0.025
r 12000_18000_M1 12000_20000_M1 0.025
r 12000_20000_M1 12000_22000_M1 0.025
r 12000_22000_M1 12000_24000_M1 0.025
r 12000_24000_M1 12000_26000_M1 0.025
r 12000_26000_M1 12000_28000_M1 0.025
r 12000_28000_M1 12000_30000_M1 0.025
r 12000_30000_M1 12000_32000_M1 0.025
r 12000_32000_M1 12000_34000_M1 0.025
r 12000_34000_M1 12000_36000_M1 0.025
r 12000_36000_M1 12000_38000_M1 0.025
r 12000_38000_M1 12000_40000_M1 0.025
r 12000_40000_M1 12000_42000_M1 0.025
r 12000_42000_M1 12000_44000_M1 0.025
r 12000_44000_M1 12000_46000_M1 0.025
r 12000_46000_M1 12000_48000_M1 0.025
r 12000_48000_M1 12000_50000_M1 0.025
r 12000_50000_M1 12000_52000_M1 0.025
r 12000_52000_M1 12000_54000_M1 0.025
r 12000_54000_M1 12000_56000_M1 0.025
r 12000_56000_M1 12000_58000_M1 0.025
r 12000_58000_M1 12000_60000_M1 0.025
r 12000_60000_M1 12000_62000_M1 0.025
r 12000_62000_M1 12000_64000_M1 0.025
r 12000_64000_M1 12000_66000_M1 0.025
r 12000_66000_M1 12000_68000_M1 0.025
r 12000_68000_M1 12000_70000_M1 0.025
r 12000_70000_M1 12000_72000_M1 0.025
r 12000_72000_M1 12000_74000_M1 0.025
r 12000_74000_M1 12000_76000_M1 0.025
r 12000_76000_M1 12000_78000_M1 0.025
r 12000_78000_M1 12000_80000_M1 0.025
r 12000_80000_M1 12000_82000_M1 0.025
r 12000_82000_M1 12000_84000_M1 0.025
r 12000_84000_M1 12000_86000_M1 0.025
r 12000_86000_M1 12000_88000_M1 0.025
r 12000_88000_M1 12000_90000_M1 0.025
r 12000_90000_M1 12000_92000_M1 0.025
r 12000_92000_M1 12000_94000_M1 0.025
r 12000_94000_M1 12000_96000_M1 0.025
r 12000_96000_M1 12000_98000_M1 0.025
r 12000_98000_M1 12000_100000_M1 0.025
r 14000_2000_M1 14000_4000_M1 0.025
r 14000_4000_M1 14000_6000_M1 0.025
r 14000_6000_M1 14000_8000_M1 0.025
r 14000_8000_M1 14000_10000_M1 0.025
r 14000_10000_M1 14000_12000_M1 0.025
r 14000_12000_M1 14000_14000_M1 0.025
r 14000_14000_M1 14000_16000_M1 0.025
r 14000_16000_M1 14000_18000_M1 0.025
r 14000_18000_M1 14000_20000_M1 0.025
r 14000_20000_M1 14000_22000_M1 0.025
r 14000_22000_M1 14000_24000_M1 0.025
r 14000_24000_M1 14000_26000_M1 0.025
r 14000_26000_M1 14000_28000_M1 0.025
r 14000_28000_M1 14000_30000_M1 0.025
r 14000_30000_M1 14000_32000_M1 0.025
r 14000_32000_M1 14000_34000_M1 0.025
r 14000_34000_M1 14000_36000_M1 0.025
r 14000_36000_M1 14000_38000_M1 0.025
r 14000_38000_M1 14000_40000_M1 0.025
r 14000_40000_M1 14000_42000_M1 0.025
r 14000_42000_M1 14000_44000_M1 0.025
r 14000_44000_M1 14000_46000_M1 0.025
r 14000_46000_M1 14000_48000_M1 0.025
r 14000_48000_M1 14000_50000_M1 0.025
r 14000_50000_M1 14000_52000_M1 0.025
r 14000_52000_M1 14000_54000_M1 0.025
r 14000_54000_M1 14000_56000_M1 0.025
r 14000_56000_M1 14000_58000_M1 0.025
r 14000_58000_M1 14000_60000_M1 0.025
r 14000_60000_M1 14000_62000_M1 0.025
r 14000_62000_M1 14000_64000_M1 0.025
r 14000_64000_M1 14000_66000_M1 0.025
r 14000_66000_M1 14000_68000_M1 0.025
r 14000_68000_M1 14000_70000_M1 0.025
r 14000_70000_M1 14000_72000_M1 0.025
r 14000_72000_M1 14000_74000_M1 0.025
r 14000_74000_M1 14000_76000_M1 0.025
r 14000_76000_M1 14000_78000_M1 0.025
r 14000_78000_M1 14000_80000_M1 0.025
r 14000_80000_M1 14000_82000_M1 0.025
r 14000_82000_M1 14000_84000_M1 0.025
r 14000_84000_M1 14000_86000_M1 0.025
r 14000_86000_M1 14000_88000_M1 0.025
r 14000_88000_M1 14000_90000_M1 0.025
r 14000_90000_M1 14000_92000_M1 0.025
r 14000_92000_M1 14000_94000_M1 0.025
r 14000_94000_M1 14000_96000_M1 0.025
r 14000_96000_M1 14000_98000_M1 0.025
r 14000_98000_M1 14000_100000_M1 0.025
r 16000_2000_M1 16000_4000_M1 0.025
r 16000_4000_M1 16000_6000_M1 0.025
r 16000_6000_M1 16000_8000_M1 0.025
r 16000_8000_M1 16000_10000_M1 0.025
r 16000_10000_M1 16000_12000_M1 0.025
r 16000_12000_M1 16000_14000_M1 0.025
r 16000_14000_M1 16000_16000_M1 0.025
r 16000_16000_M1 16000_18000_M1 0.025
r 16000_18000_M1 16000_20000_M1 0.025
r 16000_20000_M1 16000_22000_M1 0.025
r 16000_22000_M1 16000_24000_M1 0.025
r 16000_24000_M1 16000_26000_M1 0.025
r 16000_26000_M1 16000_28000_M1 0.025
r 16000_28000_M1 16000_30000_M1 0.025
r 16000_30000_M1 16000_32000_M1 0.025
r 16000_32000_M1 16000_34000_M1 0.025
r 16000_34000_M1 16000_36000_M1 0.025
r 16000_36000_M1 16000_38000_M1 0.025
r 16000_38000_M1 16000_40000_M1 0.025
r 16000_40000_M1 16000_42000_M1 0.025
r 16000_42000_M1 16000_44000_M1 0.025
r 16000_44000_M1 16000_46000_M1 0.025
r 16000_46000_M1 16000_48000_M1 0.025
r 16000_48000_M1 16000_50000_M1 0.025
r 16000_50000_M1 16000_52000_M1 0.025
r 16000_52000_M1 16000_54000_M1 0.025
r 16000_54000_M1 16000_56000_M1 0.025
r 16000_56000_M1 16000_58000_M1 0.025
r 16000_58000_M1 16000_60000_M1 0.025
r 16000_60000_M1 16000_62000_M1 0.025
r 16000_62000_M1 16000_64000_M1 0.025
r 16000_64000_M1 16000_66000_M1 0.025
r 16000_66000_M1 16000_68000_M1 0.025
r 16000_68000_M1 16000_70000_M1 0.025
r 16000_70000_M1 16000_72000_M1 0.025
r 16000_72000_M1 16000_74000_M1 0.025
r 16000_74000_M1 16000_76000_M1 0.025
r 16000_76000_M1 16000_78000_M1 0.025
r 16000_78000_M1 16000_80000_M1 0.025
r 16000_80000_M1 16000_82000_M1 0.025
r 16000_82000_M1 16000_84000_M1 0.025
r 16000_84000_M1 16000_86000_M1 0.025
r 16000_86000_M1 16000_88000_M1 0.025
r 16000_88000_M1 16000_90000_M1 0.025
r 16000_90000_M1 16000_92000_M1 0.025
r 16000_92000_M1 16000_94000_M1 0.025
r 16000_94000_M1 16000_96000_M1 0.025
r 16000_96000_M1 16000_98000_M1 0.025
r 16000_98000_M1 16000_100000_M1 0.025
r 18000_2000_M1 18000_4000_M1 0.025
r 18000_4000_M1 18000_6000_M1 0.025
r 18000_6000_M1 18000_8000_M1 0.025
r 18000_8000_M1 18000_10000_M1 0.025
r 18000_10000_M1 18000_12000_M1 0.025
r 18000_12000_M1 18000_14000_M1 0.025
r 18000_14000_M1 18000_16000_M1 0.025
r 18000_16000_M1 18000_18000_M1 0.025
r 18000_18000_M1 18000_20000_M1 0.025
r 18000_20000_M1 18000_22000_M1 0.025
r 18000_22000_M1 18000_24000_M1 0.025
r 18000_24000_M1 18000_26000_M1 0.025
r 18000_26000_M1 18000_28000_M1 0.025
r 18000_28000_M1 18000_30000_M1 0.025
r 18000_30000_M1 18000_32000_M1 0.025
r 18000_32000_M1 18000_34000_M1 0.025
r 18000_34000_M1 18000_36000_M1 0.025
r 18000_36000_M1 18000_38000_M1 0.025
r 18000_38000_M1 18000_40000_M1 0.025
r 18000_40000_M1 18000_42000_M1 0.025
r 18000_42000_M1 18000_44000_M1 0.025
r 18000_44000_M1 18000_46000_M1 0.025
r 18000_46000_M1 18000_48000_M1 0.025
r 18000_48000_M1 18000_50000_M1 0.025
r 18000_50000_M1 18000_52000_M1 0.025
r 18000_52000_M1 18000_54000_M1 0.025
r 18000_54000_M1 18000_56000_M1 0.025
r 18000_56000_M1 18000_58000_M1 0.025
r 18000_58000_M1 18000_60000_M1 0.025
r 18000_60000_M1 18000_62000_M1 0.025
r 18000_62000_M1 18000_64000_M1 0.025
r 18000_64000_M1 18000_66000_M1 0.025
r 18000_66000_M1 18000_68000_M1 0.025
r 18000_68000_M1 18000_70000_M1 0.025
r 18000_70000_M1 18000_72000_M1 0.025
r 18000_72000_M1 18000_74000_M1 0.025
r 18000_74000_M1 18000_76000_M1 0.025
r 18000_76000_M1 18000_78000_M1 0.025
r 18000_78000_M1 18000_80000_M1 0.025
r 18000_80000_M1 18000_82000_M1 0.025
r 18000_82000_M1 18000_84000_M1 0.025
r 18000_84000_M1 18000_86000_M1 0.025
r 18000_86000_M1 18000_88000_M1 0.025
r 18000_88000_M1 18000_90000_M1 0.025
r 18000_90000_M1 18000_92000_M1 0.025
r 18000_92000_M1 18000_94000_M1 0.025
r 18000_94000_M1 18000_96000_M1 0.025
r 18000_96000_M1 18000_98000_M1 0.025
r 18000_98000_M1 18000_100000_M1 0.025
r 20000_2000_M1 20000_4000_M1 0.025
r 20000_4000_M1 20000_6000_M1 0.025
r 20000_6000_M1 20000_8000_M1 0.025
r 20000_8000_M1 20000_10000_M1 0.025
r 20000_10000_M1 20000_12000_M1 0.025
r 20000_12000_M1 20000_14000_M1 0.025
r 20000_14000_M1 20000_16000_M1 0.025
r 20000_16000_M1 20000_18000_M1 0.025
r 20000_18000_M1 20000_20000_M1 0.025
r 20000_20000_M1 20000_22000_M1 0.025
r 20000_22000_M1 20000_24000_M1 0.025
r 20000_24000_M1 20000_26000_M1 0.025
r 20000_26000_M1 20000_28000_M1 0.025
r 20000_28000_M1 20000_30000_M1 0.025
r 20000_30000_M1 20000_32000_M1 0.025
r 20000_32000_M1 20000_34000_M1 0.025
r 20000_34000_M1 20000_36000_M1 0.025
r 20000_36000_M1 20000_38000_M1 0.025
r 20000_38000_M1 20000_40000_M1 0.025
r 20000_40000_M1 20000_42000_M1 0.025
r 20000_42000_M1 20000_44000_M1 0.025
r 20000_44000_M1 20000_46000_M1 0.025
r 20000_46000_M1 20000_48000_M1 0.025
r 20000_48000_M1 20000_50000_M1 0.025
r 20000_50000_M1 20000_52000_M1 0.025
r 20000_52000_M1 20000_54000_M1 0.025
r 20000_54000_M1 20000_56000_M1 0.025
r 20000_56000_M1 20000_58000_M1 0.025
r 20000_58000_M1 20000_60000_M1 0.025
r 20000_60000_M1 20000_62000_M1 0.025
r 20000_62000_M1 20000_64000_M1 0.025
r 20000_64000_M1 20000_66000_M1 0.025
r 20000_66000_M1 20000_68000_M1 0.025
r 20000_68000_M1 20000_70000_M1 0.025
r 20000_70000_M1 20000_72000_M1 0.025
r 20000_72000_M1 20000_74000_M1 0.025
r 20000_74000_M1 20000_76000_M1 0.025
r 20000_76000_M1 20000_78000_M1 0.025
r 20000_78000_M1 20000_80000_M1 0.025
r 20000_80000_M1 20000_82000_M1 0.025
r 20000_82000_M1 20000_84000_M1 0.025
r 20000_84000_M1 20000_86000_M1 0.025
r 20000_86000_M1 20000_88000_M1 0.025
r 20000_88000_M1 20000_90000_M1 0.025
r 20000_90000_M1 20000_92000_M1 0.025
r 20000_92000_M1 20000_94000_M1 0.025
r 20000_94000_M1 20000_96000_M1 0.025
r 20000_96000_M1 20000_98000_M1 0.025
r 20000_98000_M1 20000_100000_M1 0.025
r 22000_2000_M1 22000_4000_M1 0.025
r 22000_4000_M1 22000_6000_M1 0.025
r 22000_6000_M1 22000_8000_M1 0.025
r 22000_8000_M1 22000_10000_M1 0.025
r 22000_10000_M1 22000_12000_M1 0.025
r 22000_12000_M1 22000_14000_M1 0.025
r 22000_14000_M1 22000_16000_M1 0.025
r 22000_16000_M1 22000_18000_M1 0.025
r 22000_18000_M1 22000_20000_M1 0.025
r 22000_20000_M1 22000_22000_M1 0.025
r 22000_22000_M1 22000_24000_M1 0.025
r 22000_24000_M1 22000_26000_M1 0.025
r 22000_26000_M1 22000_28000_M1 0.025
r 22000_28000_M1 22000_30000_M1 0.025
r 22000_30000_M1 22000_32000_M1 0.025
r 22000_32000_M1 22000_34000_M1 0.025
r 22000_34000_M1 22000_36000_M1 0.025
r 22000_36000_M1 22000_38000_M1 0.025
r 22000_38000_M1 22000_40000_M1 0.025
r 22000_40000_M1 22000_42000_M1 0.025
r 22000_42000_M1 22000_44000_M1 0.025
r 22000_44000_M1 22000_46000_M1 0.025
r 22000_46000_M1 22000_48000_M1 0.025
r 22000_48000_M1 22000_50000_M1 0.025
r 22000_50000_M1 22000_52000_M1 0.025
r 22000_52000_M1 22000_54000_M1 0.025
r 22000_54000_M1 22000_56000_M1 0.025
r 22000_56000_M1 22000_58000_M1 0.025
r 22000_58000_M1 22000_60000_M1 0.025
r 22000_60000_M1 22000_62000_M1 0.025
r 22000_62000_M1 22000_64000_M1 0.025
r 22000_64000_M1 22000_66000_M1 0.025
r 22000_66000_M1 22000_68000_M1 0.025
r 22000_68000_M1 22000_70000_M1 0.025
r 22000_70000_M1 22000_72000_M1 0.025
r 22000_72000_M1 22000_74000_M1 0.025
r 22000_74000_M1 22000_76000_M1 0.025
r 22000_76000_M1 22000_78000_M1 0.025
r 22000_78000_M1 22000_80000_M1 0.025
r 22000_80000_M1 22000_82000_M1 0.025
r 22000_82000_M1 22000_84000_M1 0.025
r 22000_84000_M1 22000_86000_M1 0.025
r 22000_86000_M1 22000_88000_M1 0.025
r 22000_88000_M1 22000_90000_M1 0.025
r 22000_90000_M1 22000_92000_M1 0.025
r 22000_92000_M1 22000_94000_M1 0.025
r 22000_94000_M1 22000_96000_M1 0.025
r 22000_96000_M1 22000_98000_M1 0.025
r 22000_98000_M1 22000_100000_M1 0.025
r 24000_2000_M1 24000_4000_M1 0.025
r 24000_4000_M1 24000_6000_M1 0.025
r 24000_6000_M1 24000_8000_M1 0.025
r 24000_8000_M1 24000_10000_M1 0.025
r 24000_10000_M1 24000_12000_M1 0.025
r 24000_12000_M1 24000_14000_M1 0.025
r 24000_14000_M1 24000_16000_M1 0.025
r 24000_16000_M1 24000_18000_M1 0.025
r 24000_18000_M1 24000_20000_M1 0.025
r 24000_20000_M1 24000_22000_M1 0.025
r 24000_22000_M1 24000_24000_M1 0.025
r 24000_24000_M1 24000_26000_M1 0.025
r 24000_26000_M1 24000_28000_M1 0.025
r 24000_28000_M1 24000_30000_M1 0.025
r 24000_30000_M1 24000_32000_M1 0.025
r 24000_32000_M1 24000_34000_M1 0.025
r 24000_34000_M1 24000_36000_M1 0.025
r 24000_36000_M1 24000_38000_M1 0.025
r 24000_38000_M1 24000_40000_M1 0.025
r 24000_40000_M1 24000_42000_M1 0.025
r 24000_42000_M1 24000_44000_M1 0.025
r 24000_44000_M1 24000_46000_M1 0.025
r 24000_46000_M1 24000_48000_M1 0.025
r 24000_48000_M1 24000_50000_M1 0.025
r 24000_50000_M1 24000_52000_M1 0.025
r 24000_52000_M1 24000_54000_M1 0.025
r 24000_54000_M1 24000_56000_M1 0.025
r 24000_56000_M1 24000_58000_M1 0.025
r 24000_58000_M1 24000_60000_M1 0.025
r 24000_60000_M1 24000_62000_M1 0.025
r 24000_62000_M1 24000_64000_M1 0.025
r 24000_64000_M1 24000_66000_M1 0.025
r 24000_66000_M1 24000_68000_M1 0.025
r 24000_68000_M1 24000_70000_M1 0.025
r 24000_70000_M1 24000_72000_M1 0.025
r 24000_72000_M1 24000_74000_M1 0.025
r 24000_74000_M1 24000_76000_M1 0.025
r 24000_76000_M1 24000_78000_M1 0.025
r 24000_78000_M1 24000_80000_M1 0.025
r 24000_80000_M1 24000_82000_M1 0.025
r 24000_82000_M1 24000_84000_M1 0.025
r 24000_84000_M1 24000_86000_M1 0.025
r 24000_86000_M1 24000_88000_M1 0.025
r 24000_88000_M1 24000_90000_M1 0.025
r 24000_90000_M1 24000_92000_M1 0.025
r 24000_92000_M1 24000_94000_M1 0.025
r 24000_94000_M1 24000_96000_M1 0.025
r 24000_96000_M1 24000_98000_M1 0.025
r 24000_98000_M1 24000_100000_M1 0.025
r 26000_2000_M1 26000_4000_M1 0.025
r 26000_4000_M1 26000_6000_M1 0.025
r 26000_6000_M1 26000_8000_M1 0.025
r 26000_8000_M1 26000_10000_M1 0.025
r 26000_10000_M1 26000_12000_M1 0.025
r 26000_12000_M1 26000_14000_M1 0.025
r 26000_14000_M1 26000_16000_M1 0.025
r 26000_16000_M1 26000_18000_M1 0.025
r 26000_18000_M1 26000_20000_M1 0.025
r 26000_20000_M1 26000_22000_M1 0.025
r 26000_22000_M1 26000_24000_M1 0.025
r 26000_24000_M1 26000_26000_M1 0.025
r 26000_26000_M1 26000_28000_M1 0.025
r 26000_28000_M1 26000_30000_M1 0.025
r 26000_30000_M1 26000_32000_M1 0.025
r 26000_32000_M1 26000_34000_M1 0.025
r 26000_34000_M1 26000_36000_M1 0.025
r 26000_36000_M1 26000_38000_M1 0.025
r 26000_38000_M1 26000_40000_M1 0.025
r 26000_40000_M1 26000_42000_M1 0.025
r 26000_42000_M1 26000_44000_M1 0.025
r 26000_44000_M1 26000_46000_M1 0.025
r 26000_46000_M1 26000_48000_M1 0.025
r 26000_48000_M1 26000_50000_M1 0.025
r 26000_50000_M1 26000_52000_M1 0.025
r 26000_52000_M1 26000_54000_M1 0.025
r 26000_54000_M1 26000_56000_M1 0.025
r 26000_56000_M1 26000_58000_M1 0.025
r 26000_58000_M1 26000_60000_M1 0.025
r 26000_60000_M1 26000_62000_M1 0.025
r 26000_62000_M1 26000_64000_M1 0.025
r 26000_64000_M1 26000_66000_M1 0.025
r 26000_66000_M1 26000_68000_M1 0.025
r 26000_68000_M1 26000_70000_M1 0.025
r 26000_70000_M1 26000_72000_M1 0.025
r 26000_72000_M1 26000_74000_M1 0.025
r 26000_74000_M1 26000_76000_M1 0.025
r 26000_76000_M1 26000_78000_M1 0.025
r 26000_78000_M1 26000_80000_M1 0.025
r 26000_80000_M1 26000_82000_M1 0.025
r 26000_82000_M1 26000_84000_M1 0.025
r 26000_84000_M1 26000_86000_M1 0.025
r 26000_86000_M1 26000_88000_M1 0.025
r 26000_88000_M1 26000_90000_M1 0.025
r 26000_90000_M1 26000_92000_M1 0.025
r 26000_92000_M1 26000_94000_M1 0.025
r 26000_94000_M1 26000_96000_M1 0.025
r 26000_96000_M1 26000_98000_M1 0.025
r 26000_98000_M1 26000_100000_M1 0.025
r 28000_2000_M1 28000_4000_M1 0.025
r 28000_4000_M1 28000_6000_M1 0.025
r 28000_6000_M1 28000_8000_M1 0.025
r 28000_8000_M1 28000_10000_M1 0.025
r 28000_10000_M1 28000_12000_M1 0.025
r 28000_12000_M1 28000_14000_M1 0.025
r 28000_14000_M1 28000_16000_M1 0.025
r 28000_16000_M1 28000_18000_M1 0.025
r 28000_18000_M1 28000_20000_M1 0.025
r 28000_20000_M1 28000_22000_M1 0.025
r 28000_22000_M1 28000_24000_M1 0.025
r 28000_24000_M1 28000_26000_M1 0.025
r 28000_26000_M1 28000_28000_M1 0.025
r 28000_28000_M1 28000_30000_M1 0.025
r 28000_30000_M1 28000_32000_M1 0.025
r 28000_32000_M1 28000_34000_M1 0.025
r 28000_34000_M1 28000_36000_M1 0.025
r 28000_36000_M1 28000_38000_M1 0.025
r 28000_38000_M1 28000_40000_M1 0.025
r 28000_40000_M1 28000_42000_M1 0.025
r 28000_42000_M1 28000_44000_M1 0.025
r 28000_44000_M1 28000_46000_M1 0.025
r 28000_46000_M1 28000_48000_M1 0.025
r 28000_48000_M1 28000_50000_M1 0.025
r 28000_50000_M1 28000_52000_M1 0.025
r 28000_52000_M1 28000_54000_M1 0.025
r 28000_54000_M1 28000_56000_M1 0.025
r 28000_56000_M1 28000_58000_M1 0.025
r 28000_58000_M1 28000_60000_M1 0.025
r 28000_60000_M1 28000_62000_M1 0.025
r 28000_62000_M1 28000_64000_M1 0.025
r 28000_64000_M1 28000_66000_M1 0.025
r 28000_66000_M1 28000_68000_M1 0.025
r 28000_68000_M1 28000_70000_M1 0.025
r 28000_70000_M1 28000_72000_M1 0.025
r 28000_72000_M1 28000_74000_M1 0.025
r 28000_74000_M1 28000_76000_M1 0.025
r 28000_76000_M1 28000_78000_M1 0.025
r 28000_78000_M1 28000_80000_M1 0.025
r 28000_80000_M1 28000_82000_M1 0.025
r 28000_82000_M1 28000_84000_M1 0.025
r 28000_84000_M1 28000_86000_M1 0.025
r 28000_86000_M1 28000_88000_M1 0.025
r 28000_88000_M1 28000_90000_M1 0.025
r 28000_90000_M1 28000_92000_M1 0.025
r 28000_92000_M1 28000_94000_M1 0.025
r 28000_94000_M1 28000_96000_M1 0.025
r 28000_96000_M1 28000_98000_M1 0.025
r 28000_98000_M1 28000_100000_M1 0.025
r 30000_2000_M1 30000_4000_M1 0.025
r 30000_4000_M1 30000_6000_M1 0.025
r 30000_6000_M1 30000_8000_M1 0.025
r 30000_8000_M1 30000_10000_M1 0.025
r 30000_10000_M1 30000_12000_M1 0.025
r 30000_12000_M1 30000_14000_M1 0.025
r 30000_14000_M1 30000_16000_M1 0.025
r 30000_16000_M1 30000_18000_M1 0.025
r 30000_18000_M1 30000_20000_M1 0.025
r 30000_20000_M1 30000_22000_M1 0.025
r 30000_22000_M1 30000_24000_M1 0.025
r 30000_24000_M1 30000_26000_M1 0.025
r 30000_26000_M1 30000_28000_M1 0.025
r 30000_28000_M1 30000_30000_M1 0.025
r 30000_30000_M1 30000_32000_M1 0.025
r 30000_32000_M1 30000_34000_M1 0.025
r 30000_34000_M1 30000_36000_M1 0.025
r 30000_36000_M1 30000_38000_M1 0.025
r 30000_38000_M1 30000_40000_M1 0.025
r 30000_40000_M1 30000_42000_M1 0.025
r 30000_42000_M1 30000_44000_M1 0.025
r 30000_44000_M1 30000_46000_M1 0.025
r 30000_46000_M1 30000_48000_M1 0.025
r 30000_48000_M1 30000_50000_M1 0.025
r 30000_50000_M1 30000_52000_M1 0.025
r 30000_52000_M1 30000_54000_M1 0.025
r 30000_54000_M1 30000_56000_M1 0.025
r 30000_56000_M1 30000_58000_M1 0.025
r 30000_58000_M1 30000_60000_M1 0.025
r 30000_60000_M1 30000_62000_M1 0.025
r 30000_62000_M1 30000_64000_M1 0.025
r 30000_64000_M1 30000_66000_M1 0.025
r 30000_66000_M1 30000_68000_M1 0.025
r 30000_68000_M1 30000_70000_M1 0.025
r 30000_70000_M1 30000_72000_M1 0.025
r 30000_72000_M1 30000_74000_M1 0.025
r 30000_74000_M1 30000_76000_M1 0.025
r 30000_76000_M1 30000_78000_M1 0.025
r 30000_78000_M1 30000_80000_M1 0.025
r 30000_80000_M1 30000_82000_M1 0.025
r 30000_82000_M1 30000_84000_M1 0.025
r 30000_84000_M1 30000_86000_M1 0.025
r 30000_86000_M1 30000_88000_M1 0.025
r 30000_88000_M1 30000_90000_M1 0.025
r 30000_90000_M1 30000_92000_M1 0.025
r 30000_92000_M1 30000_94000_M1 0.025
r 30000_94000_M1 30000_96000_M1 0.025
r 30000_96000_M1 30000_98000_M1 0.025
r 30000_98000_M1 30000_100000_M1 0.025
r 32000_2000_M1 32000_4000_M1 0.025
r 32000_4000_M1 32000_6000_M1 0.025
r 32000_6000_M1 32000_8000_M1 0.025
r 32000_8000_M1 32000_10000_M1 0.025
r 32000_10000_M1 32000_12000_M1 0.025
r 32000_12000_M1 32000_14000_M1 0.025
r 32000_14000_M1 32000_16000_M1 0.025
r 32000_16000_M1 32000_18000_M1 0.025
r 32000_18000_M1 32000_20000_M1 0.025
r 32000_20000_M1 32000_22000_M1 0.025
r 32000_22000_M1 32000_24000_M1 0.025
r 32000_24000_M1 32000_26000_M1 0.025
r 32000_26000_M1 32000_28000_M1 0.025
r 32000_28000_M1 32000_30000_M1 0.025
r 32000_30000_M1 32000_32000_M1 0.025
r 32000_32000_M1 32000_34000_M1 0.025
r 32000_34000_M1 32000_36000_M1 0.025
r 32000_36000_M1 32000_38000_M1 0.025
r 32000_38000_M1 32000_40000_M1 0.025
r 32000_40000_M1 32000_42000_M1 0.025
r 32000_42000_M1 32000_44000_M1 0.025
r 32000_44000_M1 32000_46000_M1 0.025
r 32000_46000_M1 32000_48000_M1 0.025
r 32000_48000_M1 32000_50000_M1 0.025
r 32000_50000_M1 32000_52000_M1 0.025
r 32000_52000_M1 32000_54000_M1 0.025
r 32000_54000_M1 32000_56000_M1 0.025
r 32000_56000_M1 32000_58000_M1 0.025
r 32000_58000_M1 32000_60000_M1 0.025
r 32000_60000_M1 32000_62000_M1 0.025
r 32000_62000_M1 32000_64000_M1 0.025
r 32000_64000_M1 32000_66000_M1 0.025
r 32000_66000_M1 32000_68000_M1 0.025
r 32000_68000_M1 32000_70000_M1 0.025
r 32000_70000_M1 32000_72000_M1 0.025
r 32000_72000_M1 32000_74000_M1 0.025
r 32000_74000_M1 32000_76000_M1 0.025
r 32000_76000_M1 32000_78000_M1 0.025
r 32000_78000_M1 32000_80000_M1 0.025
r 32000_80000_M1 32000_82000_M1 0.025
r 32000_82000_M1 32000_84000_M1 0.025
r 32000_84000_M1 32000_86000_M1 0.025
r 32000_86000_M1 32000_88000_M1 0.025
r 32000_88000_M1 32000_90000_M1 0.025
r 32000_90000_M1 32000_92000_M1 0.025
r 32000_92000_M1 32000_94000_M1 0.025
r 32000_94000_M1 32000_96000_M1 0.025
r 32000_96000_M1 32000_98000_M1 0.025
r 32000_98000_M1 32000_100000_M1 0.025
r 34000_2000_M1 34000_4000_M1 0.025
r 34000_4000_M1 34000_6000_M1 0.025
r 34000_6000_M1 34000_8000_M1 0.025
r 34000_8000_M1 34000_10000_M1 0.025
r 34000_10000_M1 34000_12000_M1 0.025
r 34000_12000_M1 34000_14000_M1 0.025
r 34000_14000_M1 34000_16000_M1 0.025
r 34000_16000_M1 34000_18000_M1 0.025
r 34000_18000_M1 34000_20000_M1 0.025
r 34000_20000_M1 34000_22000_M1 0.025
r 34000_22000_M1 34000_24000_M1 0.025
r 34000_24000_M1 34000_26000_M1 0.025
r 34000_26000_M1 34000_28000_M1 0.025
r 34000_28000_M1 34000_30000_M1 0.025
r 34000_30000_M1 34000_32000_M1 0.025
r 34000_32000_M1 34000_34000_M1 0.025
r 34000_34000_M1 34000_36000_M1 0.025
r 34000_36000_M1 34000_38000_M1 0.025
r 34000_38000_M1 34000_40000_M1 0.025
r 34000_40000_M1 34000_42000_M1 0.025
r 34000_42000_M1 34000_44000_M1 0.025
r 34000_44000_M1 34000_46000_M1 0.025
r 34000_46000_M1 34000_48000_M1 0.025
r 34000_48000_M1 34000_50000_M1 0.025
r 34000_50000_M1 34000_52000_M1 0.025
r 34000_52000_M1 34000_54000_M1 0.025
r 34000_54000_M1 34000_56000_M1 0.025
r 34000_56000_M1 34000_58000_M1 0.025
r 34000_58000_M1 34000_60000_M1 0.025
r 34000_60000_M1 34000_62000_M1 0.025
r 34000_62000_M1 34000_64000_M1 0.025
r 34000_64000_M1 34000_66000_M1 0.025
r 34000_66000_M1 34000_68000_M1 0.025
r 34000_68000_M1 34000_70000_M1 0.025
r 34000_70000_M1 34000_72000_M1 0.025
r 34000_72000_M1 34000_74000_M1 0.025
r 34000_74000_M1 34000_76000_M1 0.025
r 34000_76000_M1 34000_78000_M1 0.025
r 34000_78000_M1 34000_80000_M1 0.025
r 34000_80000_M1 34000_82000_M1 0.025
r 34000_82000_M1 34000_84000_M1 0.025
r 34000_84000_M1 34000_86000_M1 0.025
r 34000_86000_M1 34000_88000_M1 0.025
r 34000_88000_M1 34000_90000_M1 0.025
r 34000_90000_M1 34000_92000_M1 0.025
r 34000_92000_M1 34000_94000_M1 0.025
r 34000_94000_M1 34000_96000_M1 0.025
r 34000_96000_M1 34000_98000_M1 0.025
r 34000_98000_M1 34000_100000_M1 0.025
r 36000_2000_M1 36000_4000_M1 0.025
r 36000_4000_M1 36000_6000_M1 0.025
r 36000_6000_M1 36000_8000_M1 0.025
r 36000_8000_M1 36000_10000_M1 0.025
r 36000_10000_M1 36000_12000_M1 0.025
r 36000_12000_M1 36000_14000_M1 0.025
r 36000_14000_M1 36000_16000_M1 0.025
r 36000_16000_M1 36000_18000_M1 0.025
r 36000_18000_M1 36000_20000_M1 0.025
r 36000_20000_M1 36000_22000_M1 0.025
r 36000_22000_M1 36000_24000_M1 0.025
r 36000_24000_M1 36000_26000_M1 0.025
r 36000_26000_M1 36000_28000_M1 0.025
r 36000_28000_M1 36000_30000_M1 0.025
r 36000_30000_M1 36000_32000_M1 0.025
r 36000_32000_M1 36000_34000_M1 0.025
r 36000_34000_M1 36000_36000_M1 0.025
r 36000_36000_M1 36000_38000_M1 0.025
r 36000_38000_M1 36000_40000_M1 0.025
r 36000_40000_M1 36000_42000_M1 0.025
r 36000_42000_M1 36000_44000_M1 0.025
r 36000_44000_M1 36000_46000_M1 0.025
r 36000_46000_M1 36000_48000_M1 0.025
r 36000_48000_M1 36000_50000_M1 0.025
r 36000_50000_M1 36000_52000_M1 0.025
r 36000_52000_M1 36000_54000_M1 0.025
r 36000_54000_M1 36000_56000_M1 0.025
r 36000_56000_M1 36000_58000_M1 0.025
r 36000_58000_M1 36000_60000_M1 0.025
r 36000_60000_M1 36000_62000_M1 0.025
r 36000_62000_M1 36000_64000_M1 0.025
r 36000_64000_M1 36000_66000_M1 0.025
r 36000_66000_M1 36000_68000_M1 0.025
r 36000_68000_M1 36000_70000_M1 0.025
r 36000_70000_M1 36000_72000_M1 0.025
r 36000_72000_M1 36000_74000_M1 0.025
r 36000_74000_M1 36000_76000_M1 0.025
r 36000_76000_M1 36000_78000_M1 0.025
r 36000_78000_M1 36000_80000_M1 0.025
r 36000_80000_M1 36000_82000_M1 0.025
r 36000_82000_M1 36000_84000_M1 0.025
r 36000_84000_M1 36000_86000_M1 0.025
r 36000_86000_M1 36000_88000_M1 0.025
r 36000_88000_M1 36000_90000_M1 0.025
r 36000_90000_M1 36000_92000_M1 0.025
r 36000_92000_M1 36000_94000_M1 0.025
r 36000_94000_M1 36000_96000_M1 0.025
r 36000_96000_M1 36000_98000_M1 0.025
r 36000_98000_M1 36000_100000_M1 0.025
r 38000_2000_M1 38000_4000_M1 0.025
r 38000_4000_M1 38000_6000_M1 0.025
r 38000_6000_M1 38000_8000_M1 0.025
r 38000_8000_M1 38000_10000_M1 0.025
r 38000_10000_M1 38000_12000_M1 0.025
r 38000_12000_M1 38000_14000_M1 0.025
r 38000_14000_M1 38000_16000_M1 0.025
r 38000_16000_M1 38000_18000_M1 0.025
r 38000_18000_M1 38000_20000_M1 0.025
r 38000_20000_M1 38000_22000_M1 0.025
r 38000_22000_M1 38000_24000_M1 0.025
r 38000_24000_M1 38000_26000_M1 0.025
r 38000_26000_M1 38000_28000_M1 0.025
r 38000_28000_M1 38000_30000_M1 0.025
r 38000_30000_M1 38000_32000_M1 0.025
r 38000_32000_M1 38000_34000_M1 0.025
r 38000_34000_M1 38000_36000_M1 0.025
r 38000_36000_M1 38000_38000_M1 0.025
r 38000_38000_M1 38000_40000_M1 0.025
r 38000_40000_M1 38000_42000_M1 0.025
r 38000_42000_M1 38000_44000_M1 0.025
r 38000_44000_M1 38000_46000_M1 0.025
r 38000_46000_M1 38000_48000_M1 0.025
r 38000_48000_M1 38000_50000_M1 0.025
r 38000_50000_M1 38000_52000_M1 0.025
r 38000_52000_M1 38000_54000_M1 0.025
r 38000_54000_M1 38000_56000_M1 0.025
r 38000_56000_M1 38000_58000_M1 0.025
r 38000_58000_M1 38000_60000_M1 0.025
r 38000_60000_M1 38000_62000_M1 0.025
r 38000_62000_M1 38000_64000_M1 0.025
r 38000_64000_M1 38000_66000_M1 0.025
r 38000_66000_M1 38000_68000_M1 0.025
r 38000_68000_M1 38000_70000_M1 0.025
r 38000_70000_M1 38000_72000_M1 0.025
r 38000_72000_M1 38000_74000_M1 0.025
r 38000_74000_M1 38000_76000_M1 0.025
r 38000_76000_M1 38000_78000_M1 0.025
r 38000_78000_M1 38000_80000_M1 0.025
r 38000_80000_M1 38000_82000_M1 0.025
r 38000_82000_M1 38000_84000_M1 0.025
r 38000_84000_M1 38000_86000_M1 0.025
r 38000_86000_M1 38000_88000_M1 0.025
r 38000_88000_M1 38000_90000_M1 0.025
r 38000_90000_M1 38000_92000_M1 0.025
r 38000_92000_M1 38000_94000_M1 0.025
r 38000_94000_M1 38000_96000_M1 0.025
r 38000_96000_M1 38000_98000_M1 0.025
r 38000_98000_M1 38000_100000_M1 0.025
r 40000_2000_M1 40000_4000_M1 0.025
r 40000_4000_M1 40000_6000_M1 0.025
r 40000_6000_M1 40000_8000_M1 0.025
r 40000_8000_M1 40000_10000_M1 0.025
r 40000_10000_M1 40000_12000_M1 0.025
r 40000_12000_M1 40000_14000_M1 0.025
r 40000_14000_M1 40000_16000_M1 0.025
r 40000_16000_M1 40000_18000_M1 0.025
r 40000_18000_M1 40000_20000_M1 0.025
r 40000_20000_M1 40000_22000_M1 0.025
r 40000_22000_M1 40000_24000_M1 0.025
r 40000_24000_M1 40000_26000_M1 0.025
r 40000_26000_M1 40000_28000_M1 0.025
r 40000_28000_M1 40000_30000_M1 0.025
r 40000_30000_M1 40000_32000_M1 0.025
r 40000_32000_M1 40000_34000_M1 0.025
r 40000_34000_M1 40000_36000_M1 0.025
r 40000_36000_M1 40000_38000_M1 0.025
r 40000_38000_M1 40000_40000_M1 0.025
r 40000_40000_M1 40000_42000_M1 0.025
r 40000_42000_M1 40000_44000_M1 0.025
r 40000_44000_M1 40000_46000_M1 0.025
r 40000_46000_M1 40000_48000_M1 0.025
r 40000_48000_M1 40000_50000_M1 0.025
r 40000_50000_M1 40000_52000_M1 0.025
r 40000_52000_M1 40000_54000_M1 0.025
r 40000_54000_M1 40000_56000_M1 0.025
r 40000_56000_M1 40000_58000_M1 0.025
r 40000_58000_M1 40000_60000_M1 0.025
r 40000_60000_M1 40000_62000_M1 0.025
r 40000_62000_M1 40000_64000_M1 0.025
r 40000_64000_M1 40000_66000_M1 0.025
r 40000_66000_M1 40000_68000_M1 0.025
r 40000_68000_M1 40000_70000_M1 0.025
r 40000_70000_M1 40000_72000_M1 0.025
r 40000_72000_M1 40000_74000_M1 0.025
r 40000_74000_M1 40000_76000_M1 0.025
r 40000_76000_M1 40000_78000_M1 0.025
r 40000_78000_M1 40000_80000_M1 0.025
r 40000_80000_M1 40000_82000_M1 0.025
r 40000_82000_M1 40000_84000_M1 0.025
r 40000_84000_M1 40000_86000_M1 0.025
r 40000_86000_M1 40000_88000_M1 0.025
r 40000_88000_M1 40000_90000_M1 0.025
r 40000_90000_M1 40000_92000_M1 0.025
r 40000_92000_M1 40000_94000_M1 0.025
r 40000_94000_M1 40000_96000_M1 0.025
r 40000_96000_M1 40000_98000_M1 0.025
r 40000_98000_M1 40000_100000_M1 0.025
r 42000_2000_M1 42000_4000_M1 0.025
r 42000_4000_M1 42000_6000_M1 0.025
r 42000_6000_M1 42000_8000_M1 0.025
r 42000_8000_M1 42000_10000_M1 0.025
r 42000_10000_M1 42000_12000_M1 0.025
r 42000_12000_M1 42000_14000_M1 0.025
r 42000_14000_M1 42000_16000_M1 0.025
r 42000_16000_M1 42000_18000_M1 0.025
r 42000_18000_M1 42000_20000_M1 0.025
r 42000_20000_M1 42000_22000_M1 0.025
r 42000_22000_M1 42000_24000_M1 0.025
r 42000_24000_M1 42000_26000_M1 0.025
r 42000_26000_M1 42000_28000_M1 0.025
r 42000_28000_M1 42000_30000_M1 0.025
r 42000_30000_M1 42000_32000_M1 0.025
r 42000_32000_M1 42000_34000_M1 0.025
r 42000_34000_M1 42000_36000_M1 0.025
r 42000_36000_M1 42000_38000_M1 0.025
r 42000_38000_M1 42000_40000_M1 0.025
r 42000_40000_M1 42000_42000_M1 0.025
r 42000_42000_M1 42000_44000_M1 0.025
r 42000_44000_M1 42000_46000_M1 0.025
r 42000_46000_M1 42000_48000_M1 0.025
r 42000_48000_M1 42000_50000_M1 0.025
r 42000_50000_M1 42000_52000_M1 0.025
r 42000_52000_M1 42000_54000_M1 0.025
r 42000_54000_M1 42000_56000_M1 0.025
r 42000_56000_M1 42000_58000_M1 0.025
r 42000_58000_M1 42000_60000_M1 0.025
r 42000_60000_M1 42000_62000_M1 0.025
r 42000_62000_M1 42000_64000_M1 0.025
r 42000_64000_M1 42000_66000_M1 0.025
r 42000_66000_M1 42000_68000_M1 0.025
r 42000_68000_M1 42000_70000_M1 0.025
r 42000_70000_M1 42000_72000_M1 0.025
r 42000_72000_M1 42000_74000_M1 0.025
r 42000_74000_M1 42000_76000_M1 0.025
r 42000_76000_M1 42000_78000_M1 0.025
r 42000_78000_M1 42000_80000_M1 0.025
r 42000_80000_M1 42000_82000_M1 0.025
r 42000_82000_M1 42000_84000_M1 0.025
r 42000_84000_M1 42000_86000_M1 0.025
r 42000_86000_M1 42000_88000_M1 0.025
r 42000_88000_M1 42000_90000_M1 0.025
r 42000_90000_M1 42000_92000_M1 0.025
r 42000_92000_M1 42000_94000_M1 0.025
r 42000_94000_M1 42000_96000_M1 0.025
r 42000_96000_M1 42000_98000_M1 0.025
r 42000_98000_M1 42000_100000_M1 0.025
r 44000_2000_M1 44000_4000_M1 0.025
r 44000_4000_M1 44000_6000_M1 0.025
r 44000_6000_M1 44000_8000_M1 0.025
r 44000_8000_M1 44000_10000_M1 0.025
r 44000_10000_M1 44000_12000_M1 0.025
r 44000_12000_M1 44000_14000_M1 0.025
r 44000_14000_M1 44000_16000_M1 0.025
r 44000_16000_M1 44000_18000_M1 0.025
r 44000_18000_M1 44000_20000_M1 0.025
r 44000_20000_M1 44000_22000_M1 0.025
r 44000_22000_M1 44000_24000_M1 0.025
r 44000_24000_M1 44000_26000_M1 0.025
r 44000_26000_M1 44000_28000_M1 0.025
r 44000_28000_M1 44000_30000_M1 0.025
r 44000_30000_M1 44000_32000_M1 0.025
r 44000_32000_M1 44000_34000_M1 0.025
r 44000_34000_M1 44000_36000_M1 0.025
r 44000_36000_M1 44000_38000_M1 0.025
r 44000_38000_M1 44000_40000_M1 0.025
r 44000_40000_M1 44000_42000_M1 0.025
r 44000_42000_M1 44000_44000_M1 0.025
r 44000_44000_M1 44000_46000_M1 0.025
r 44000_46000_M1 44000_48000_M1 0.025
r 44000_48000_M1 44000_50000_M1 0.025
r 44000_50000_M1 44000_52000_M1 0.025
r 44000_52000_M1 44000_54000_M1 0.025
r 44000_54000_M1 44000_56000_M1 0.025
r 44000_56000_M1 44000_58000_M1 0.025
r 44000_58000_M1 44000_60000_M1 0.025
r 44000_60000_M1 44000_62000_M1 0.025
r 44000_62000_M1 44000_64000_M1 0.025
r 44000_64000_M1 44000_66000_M1 0.025
r 44000_66000_M1 44000_68000_M1 0.025
r 44000_68000_M1 44000_70000_M1 0.025
r 44000_70000_M1 44000_72000_M1 0.025
r 44000_72000_M1 44000_74000_M1 0.025
r 44000_74000_M1 44000_76000_M1 0.025
r 44000_76000_M1 44000_78000_M1 0.025
r 44000_78000_M1 44000_80000_M1 0.025
r 44000_80000_M1 44000_82000_M1 0.025
r 44000_82000_M1 44000_84000_M1 0.025
r 44000_84000_M1 44000_86000_M1 0.025
r 44000_86000_M1 44000_88000_M1 0.025
r 44000_88000_M1 44000_90000_M1 0.025
r 44000_90000_M1 44000_92000_M1 0.025
r 44000_92000_M1 44000_94000_M1 0.025
r 44000_94000_M1 44000_96000_M1 0.025
r 44000_96000_M1 44000_98000_M1 0.025
r 44000_98000_M1 44000_100000_M1 0.025
r 46000_2000_M1 46000_4000_M1 0.025
r 46000_4000_M1 46000_6000_M1 0.025
r 46000_6000_M1 46000_8000_M1 0.025
r 46000_8000_M1 46000_10000_M1 0.025
r 46000_10000_M1 46000_12000_M1 0.025
r 46000_12000_M1 46000_14000_M1 0.025
r 46000_14000_M1 46000_16000_M1 0.025
r 46000_16000_M1 46000_18000_M1 0.025
r 46000_18000_M1 46000_20000_M1 0.025
r 46000_20000_M1 46000_22000_M1 0.025
r 46000_22000_M1 46000_24000_M1 0.025
r 46000_24000_M1 46000_26000_M1 0.025
r 46000_26000_M1 46000_28000_M1 0.025
r 46000_28000_M1 46000_30000_M1 0.025
r 46000_30000_M1 46000_32000_M1 0.025
r 46000_32000_M1 46000_34000_M1 0.025
r 46000_34000_M1 46000_36000_M1 0.025
r 46000_36000_M1 46000_38000_M1 0.025
r 46000_38000_M1 46000_40000_M1 0.025
r 46000_40000_M1 46000_42000_M1 0.025
r 46000_42000_M1 46000_44000_M1 0.025
r 46000_44000_M1 46000_46000_M1 0.025
r 46000_46000_M1 46000_48000_M1 0.025
r 46000_48000_M1 46000_50000_M1 0.025
r 46000_50000_M1 46000_52000_M1 0.025
r 46000_52000_M1 46000_54000_M1 0.025
r 46000_54000_M1 46000_56000_M1 0.025
r 46000_56000_M1 46000_58000_M1 0.025
r 46000_58000_M1 46000_60000_M1 0.025
r 46000_60000_M1 46000_62000_M1 0.025
r 46000_62000_M1 46000_64000_M1 0.025
r 46000_64000_M1 46000_66000_M1 0.025
r 46000_66000_M1 46000_68000_M1 0.025
r 46000_68000_M1 46000_70000_M1 0.025
r 46000_70000_M1 46000_72000_M1 0.025
r 46000_72000_M1 46000_74000_M1 0.025
r 46000_74000_M1 46000_76000_M1 0.025
r 46000_76000_M1 46000_78000_M1 0.025
r 46000_78000_M1 46000_80000_M1 0.025
r 46000_80000_M1 46000_82000_M1 0.025
r 46000_82000_M1 46000_84000_M1 0.025
r 46000_84000_M1 46000_86000_M1 0.025
r 46000_86000_M1 46000_88000_M1 0.025
r 46000_88000_M1 46000_90000_M1 0.025
r 46000_90000_M1 46000_92000_M1 0.025
r 46000_92000_M1 46000_94000_M1 0.025
r 46000_94000_M1 46000_96000_M1 0.025
r 46000_96000_M1 46000_98000_M1 0.025
r 46000_98000_M1 46000_100000_M1 0.025
r 48000_2000_M1 48000_4000_M1 0.025
r 48000_4000_M1 48000_6000_M1 0.025
r 48000_6000_M1 48000_8000_M1 0.025
r 48000_8000_M1 48000_10000_M1 0.025
r 48000_10000_M1 48000_12000_M1 0.025
r 48000_12000_M1 48000_14000_M1 0.025
r 48000_14000_M1 48000_16000_M1 0.025
r 48000_16000_M1 48000_18000_M1 0.025
r 48000_18000_M1 48000_20000_M1 0.025
r 48000_20000_M1 48000_22000_M1 0.025
r 48000_22000_M1 48000_24000_M1 0.025
r 48000_24000_M1 48000_26000_M1 0.025
r 48000_26000_M1 48000_28000_M1 0.025
r 48000_28000_M1 48000_30000_M1 0.025
r 48000_30000_M1 48000_32000_M1 0.025
r 48000_32000_M1 48000_34000_M1 0.025
r 48000_34000_M1 48000_36000_M1 0.025
r 48000_36000_M1 48000_38000_M1 0.025
r 48000_38000_M1 48000_40000_M1 0.025
r 48000_40000_M1 48000_42000_M1 0.025
r 48000_42000_M1 48000_44000_M1 0.025
r 48000_44000_M1 48000_46000_M1 0.025
r 48000_46000_M1 48000_48000_M1 0.025
r 48000_48000_M1 48000_50000_M1 0.025
r 48000_50000_M1 48000_52000_M1 0.025
r 48000_52000_M1 48000_54000_M1 0.025
r 48000_54000_M1 48000_56000_M1 0.025
r 48000_56000_M1 48000_58000_M1 0.025
r 48000_58000_M1 48000_60000_M1 0.025
r 48000_60000_M1 48000_62000_M1 0.025
r 48000_62000_M1 48000_64000_M1 0.025
r 48000_64000_M1 48000_66000_M1 0.025
r 48000_66000_M1 48000_68000_M1 0.025
r 48000_68000_M1 48000_70000_M1 0.025
r 48000_70000_M1 48000_72000_M1 0.025
r 48000_72000_M1 48000_74000_M1 0.025
r 48000_74000_M1 48000_76000_M1 0.025
r 48000_76000_M1 48000_78000_M1 0.025
r 48000_78000_M1 48000_80000_M1 0.025
r 48000_80000_M1 48000_82000_M1 0.025
r 48000_82000_M1 48000_84000_M1 0.025
r 48000_84000_M1 48000_86000_M1 0.025
r 48000_86000_M1 48000_88000_M1 0.025
r 48000_88000_M1 48000_90000_M1 0.025
r 48000_90000_M1 48000_92000_M1 0.025
r 48000_92000_M1 48000_94000_M1 0.025
r 48000_94000_M1 48000_96000_M1 0.025
r 48000_96000_M1 48000_98000_M1 0.025
r 48000_98000_M1 48000_100000_M1 0.025
r 50000_2000_M1 50000_4000_M1 0.025
r 50000_4000_M1 50000_6000_M1 0.025
r 50000_6000_M1 50000_8000_M1 0.025
r 50000_8000_M1 50000_10000_M1 0.025
r 50000_10000_M1 50000_12000_M1 0.025
r 50000_12000_M1 50000_14000_M1 0.025
r 50000_14000_M1 50000_16000_M1 0.025
r 50000_16000_M1 50000_18000_M1 0.025
r 50000_18000_M1 50000_20000_M1 0.025
r 50000_20000_M1 50000_22000_M1 0.025
r 50000_22000_M1 50000_24000_M1 0.025
r 50000_24000_M1 50000_26000_M1 0.025
r 50000_26000_M1 50000_28000_M1 0.025
r 50000_28000_M1 50000_30000_M1 0.025
r 50000_30000_M1 50000_32000_M1 0.025
r 50000_32000_M1 50000_34000_M1 0.025
r 50000_34000_M1 50000_36000_M1 0.025
r 50000_36000_M1 50000_38000_M1 0.025
r 50000_38000_M1 50000_40000_M1 0.025
r 50000_40000_M1 50000_42000_M1 0.025
r 50000_42000_M1 50000_44000_M1 0.025
r 50000_44000_M1 50000_46000_M1 0.025
r 50000_46000_M1 50000_48000_M1 0.025
r 50000_48000_M1 50000_50000_M1 0.025
r 50000_50000_M1 50000_52000_M1 0.025
r 50000_52000_M1 50000_54000_M1 0.025
r 50000_54000_M1 50000_56000_M1 0.025
r 50000_56000_M1 50000_58000_M1 0.025
r 50000_58000_M1 50000_60000_M1 0.025
r 50000_60000_M1 50000_62000_M1 0.025
r 50000_62000_M1 50000_64000_M1 0.025
r 50000_64000_M1 50000_66000_M1 0.025
r 50000_66000_M1 50000_68000_M1 0.025
r 50000_68000_M1 50000_70000_M1 0.025
r 50000_70000_M1 50000_72000_M1 0.025
r 50000_72000_M1 50000_74000_M1 0.025
r 50000_74000_M1 50000_76000_M1 0.025
r 50000_76000_M1 50000_78000_M1 0.025
r 50000_78000_M1 50000_80000_M1 0.025
r 50000_80000_M1 50000_82000_M1 0.025
r 50000_82000_M1 50000_84000_M1 0.025
r 50000_84000_M1 50000_86000_M1 0.025
r 50000_86000_M1 50000_88000_M1 0.025
r 50000_88000_M1 50000_90000_M1 0.025
r 50000_90000_M1 50000_92000_M1 0.025
r 50000_92000_M1 50000_94000_M1 0.025
r 50000_94000_M1 50000_96000_M1 0.025
r 50000_96000_M1 50000_98000_M1 0.025
r 50000_98000_M1 50000_100000_M1 0.025
r 52000_2000_M1 52000_4000_M1 0.025
r 52000_4000_M1 52000_6000_M1 0.025
r 52000_6000_M1 52000_8000_M1 0.025
r 52000_8000_M1 52000_10000_M1 0.025
r 52000_10000_M1 52000_12000_M1 0.025
r 52000_12000_M1 52000_14000_M1 0.025
r 52000_14000_M1 52000_16000_M1 0.025
r 52000_16000_M1 52000_18000_M1 0.025
r 52000_18000_M1 52000_20000_M1 0.025
r 52000_20000_M1 52000_22000_M1 0.025
r 52000_22000_M1 52000_24000_M1 0.025
r 52000_24000_M1 52000_26000_M1 0.025
r 52000_26000_M1 52000_28000_M1 0.025
r 52000_28000_M1 52000_30000_M1 0.025
r 52000_30000_M1 52000_32000_M1 0.025
r 52000_32000_M1 52000_34000_M1 0.025
r 52000_34000_M1 52000_36000_M1 0.025
r 52000_36000_M1 52000_38000_M1 0.025
r 52000_38000_M1 52000_40000_M1 0.025
r 52000_40000_M1 52000_42000_M1 0.025
r 52000_42000_M1 52000_44000_M1 0.025
r 52000_44000_M1 52000_46000_M1 0.025
r 52000_46000_M1 52000_48000_M1 0.025
r 52000_48000_M1 52000_50000_M1 0.025
r 52000_50000_M1 52000_52000_M1 0.025
r 52000_52000_M1 52000_54000_M1 0.025
r 52000_54000_M1 52000_56000_M1 0.025
r 52000_56000_M1 52000_58000_M1 0.025
r 52000_58000_M1 52000_60000_M1 0.025
r 52000_60000_M1 52000_62000_M1 0.025
r 52000_62000_M1 52000_64000_M1 0.025
r 52000_64000_M1 52000_66000_M1 0.025
r 52000_66000_M1 52000_68000_M1 0.025
r 52000_68000_M1 52000_70000_M1 0.025
r 52000_70000_M1 52000_72000_M1 0.025
r 52000_72000_M1 52000_74000_M1 0.025
r 52000_74000_M1 52000_76000_M1 0.025
r 52000_76000_M1 52000_78000_M1 0.025
r 52000_78000_M1 52000_80000_M1 0.025
r 52000_80000_M1 52000_82000_M1 0.025
r 52000_82000_M1 52000_84000_M1 0.025
r 52000_84000_M1 52000_86000_M1 0.025
r 52000_86000_M1 52000_88000_M1 0.025
r 52000_88000_M1 52000_90000_M1 0.025
r 52000_90000_M1 52000_92000_M1 0.025
r 52000_92000_M1 52000_94000_M1 0.025
r 52000_94000_M1 52000_96000_M1 0.025
r 52000_96000_M1 52000_98000_M1 0.025
r 52000_98000_M1 52000_100000_M1 0.025
r 54000_2000_M1 54000_4000_M1 0.025
r 54000_4000_M1 54000_6000_M1 0.025
r 54000_6000_M1 54000_8000_M1 0.025
r 54000_8000_M1 54000_10000_M1 0.025
r 54000_10000_M1 54000_12000_M1 0.025
r 54000_12000_M1 54000_14000_M1 0.025
r 54000_14000_M1 54000_16000_M1 0.025
r 54000_16000_M1 54000_18000_M1 0.025
r 54000_18000_M1 54000_20000_M1 0.025
r 54000_20000_M1 54000_22000_M1 0.025
r 54000_22000_M1 54000_24000_M1 0.025
r 54000_24000_M1 54000_26000_M1 0.025
r 54000_26000_M1 54000_28000_M1 0.025
r 54000_28000_M1 54000_30000_M1 0.025
r 54000_30000_M1 54000_32000_M1 0.025
r 54000_32000_M1 54000_34000_M1 0.025
r 54000_34000_M1 54000_36000_M1 0.025
r 54000_36000_M1 54000_38000_M1 0.025
r 54000_38000_M1 54000_40000_M1 0.025
r 54000_40000_M1 54000_42000_M1 0.025
r 54000_42000_M1 54000_44000_M1 0.025
r 54000_44000_M1 54000_46000_M1 0.025
r 54000_46000_M1 54000_48000_M1 0.025
r 54000_48000_M1 54000_50000_M1 0.025
r 54000_50000_M1 54000_52000_M1 0.025
r 54000_52000_M1 54000_54000_M1 0.025
r 54000_54000_M1 54000_56000_M1 0.025
r 54000_56000_M1 54000_58000_M1 0.025
r 54000_58000_M1 54000_60000_M1 0.025
r 54000_60000_M1 54000_62000_M1 0.025
r 54000_62000_M1 54000_64000_M1 0.025
r 54000_64000_M1 54000_66000_M1 0.025
r 54000_66000_M1 54000_68000_M1 0.025
r 54000_68000_M1 54000_70000_M1 0.025
r 54000_70000_M1 54000_72000_M1 0.025
r 54000_72000_M1 54000_74000_M1 0.025
r 54000_74000_M1 54000_76000_M1 0.025
r 54000_76000_M1 54000_78000_M1 0.025
r 54000_78000_M1 54000_80000_M1 0.025
r 54000_80000_M1 54000_82000_M1 0.025
r 54000_82000_M1 54000_84000_M1 0.025
r 54000_84000_M1 54000_86000_M1 0.025
r 54000_86000_M1 54000_88000_M1 0.025
r 54000_88000_M1 54000_90000_M1 0.025
r 54000_90000_M1 54000_92000_M1 0.025
r 54000_92000_M1 54000_94000_M1 0.025
r 54000_94000_M1 54000_96000_M1 0.025
r 54000_96000_M1 54000_98000_M1 0.025
r 54000_98000_M1 54000_100000_M1 0.025
r 56000_2000_M1 56000_4000_M1 0.025
r 56000_4000_M1 56000_6000_M1 0.025
r 56000_6000_M1 56000_8000_M1 0.025
r 56000_8000_M1 56000_10000_M1 0.025
r 56000_10000_M1 56000_12000_M1 0.025
r 56000_12000_M1 56000_14000_M1 0.025
r 56000_14000_M1 56000_16000_M1 0.025
r 56000_16000_M1 56000_18000_M1 0.025
r 56000_18000_M1 56000_20000_M1 0.025
r 56000_20000_M1 56000_22000_M1 0.025
r 56000_22000_M1 56000_24000_M1 0.025
r 56000_24000_M1 56000_26000_M1 0.025
r 56000_26000_M1 56000_28000_M1 0.025
r 56000_28000_M1 56000_30000_M1 0.025
r 56000_30000_M1 56000_32000_M1 0.025
r 56000_32000_M1 56000_34000_M1 0.025
r 56000_34000_M1 56000_36000_M1 0.025
r 56000_36000_M1 56000_38000_M1 0.025
r 56000_38000_M1 56000_40000_M1 0.025
r 56000_40000_M1 56000_42000_M1 0.025
r 56000_42000_M1 56000_44000_M1 0.025
r 56000_44000_M1 56000_46000_M1 0.025
r 56000_46000_M1 56000_48000_M1 0.025
r 56000_48000_M1 56000_50000_M1 0.025
r 56000_50000_M1 56000_52000_M1 0.025
r 56000_52000_M1 56000_54000_M1 0.025
r 56000_54000_M1 56000_56000_M1 0.025
r 56000_56000_M1 56000_58000_M1 0.025
r 56000_58000_M1 56000_60000_M1 0.025
r 56000_60000_M1 56000_62000_M1 0.025
r 56000_62000_M1 56000_64000_M1 0.025
r 56000_64000_M1 56000_66000_M1 0.025
r 56000_66000_M1 56000_68000_M1 0.025
r 56000_68000_M1 56000_70000_M1 0.025
r 56000_70000_M1 56000_72000_M1 0.025
r 56000_72000_M1 56000_74000_M1 0.025
r 56000_74000_M1 56000_76000_M1 0.025
r 56000_76000_M1 56000_78000_M1 0.025
r 56000_78000_M1 56000_80000_M1 0.025
r 56000_80000_M1 56000_82000_M1 0.025
r 56000_82000_M1 56000_84000_M1 0.025
r 56000_84000_M1 56000_86000_M1 0.025
r 56000_86000_M1 56000_88000_M1 0.025
r 56000_88000_M1 56000_90000_M1 0.025
r 56000_90000_M1 56000_92000_M1 0.025
r 56000_92000_M1 56000_94000_M1 0.025
r 56000_94000_M1 56000_96000_M1 0.025
r 56000_96000_M1 56000_98000_M1 0.025
r 56000_98000_M1 56000_100000_M1 0.025
r 58000_2000_M1 58000_4000_M1 0.025
r 58000_4000_M1 58000_6000_M1 0.025
r 58000_6000_M1 58000_8000_M1 0.025
r 58000_8000_M1 58000_10000_M1 0.025
r 58000_10000_M1 58000_12000_M1 0.025
r 58000_12000_M1 58000_14000_M1 0.025
r 58000_14000_M1 58000_16000_M1 0.025
r 58000_16000_M1 58000_18000_M1 0.025
r 58000_18000_M1 58000_20000_M1 0.025
r 58000_20000_M1 58000_22000_M1 0.025
r 58000_22000_M1 58000_24000_M1 0.025
r 58000_24000_M1 58000_26000_M1 0.025
r 58000_26000_M1 58000_28000_M1 0.025
r 58000_28000_M1 58000_30000_M1 0.025
r 58000_30000_M1 58000_32000_M1 0.025
r 58000_32000_M1 58000_34000_M1 0.025
r 58000_34000_M1 58000_36000_M1 0.025
r 58000_36000_M1 58000_38000_M1 0.025
r 58000_38000_M1 58000_40000_M1 0.025
r 58000_40000_M1 58000_42000_M1 0.025
r 58000_42000_M1 58000_44000_M1 0.025
r 58000_44000_M1 58000_46000_M1 0.025
r 58000_46000_M1 58000_48000_M1 0.025
r 58000_48000_M1 58000_50000_M1 0.025
r 58000_50000_M1 58000_52000_M1 0.025
r 58000_52000_M1 58000_54000_M1 0.025
r 58000_54000_M1 58000_56000_M1 0.025
r 58000_56000_M1 58000_58000_M1 0.025
r 58000_58000_M1 58000_60000_M1 0.025
r 58000_60000_M1 58000_62000_M1 0.025
r 58000_62000_M1 58000_64000_M1 0.025
r 58000_64000_M1 58000_66000_M1 0.025
r 58000_66000_M1 58000_68000_M1 0.025
r 58000_68000_M1 58000_70000_M1 0.025
r 58000_70000_M1 58000_72000_M1 0.025
r 58000_72000_M1 58000_74000_M1 0.025
r 58000_74000_M1 58000_76000_M1 0.025
r 58000_76000_M1 58000_78000_M1 0.025
r 58000_78000_M1 58000_80000_M1 0.025
r 58000_80000_M1 58000_82000_M1 0.025
r 58000_82000_M1 58000_84000_M1 0.025
r 58000_84000_M1 58000_86000_M1 0.025
r 58000_86000_M1 58000_88000_M1 0.025
r 58000_88000_M1 58000_90000_M1 0.025
r 58000_90000_M1 58000_92000_M1 0.025
r 58000_92000_M1 58000_94000_M1 0.025
r 58000_94000_M1 58000_96000_M1 0.025
r 58000_96000_M1 58000_98000_M1 0.025
r 58000_98000_M1 58000_100000_M1 0.025
r 60000_2000_M1 60000_4000_M1 0.025
r 60000_4000_M1 60000_6000_M1 0.025
r 60000_6000_M1 60000_8000_M1 0.025
r 60000_8000_M1 60000_10000_M1 0.025
r 60000_10000_M1 60000_12000_M1 0.025
r 60000_12000_M1 60000_14000_M1 0.025
r 60000_14000_M1 60000_16000_M1 0.025
r 60000_16000_M1 60000_18000_M1 0.025
r 60000_18000_M1 60000_20000_M1 0.025
r 60000_20000_M1 60000_22000_M1 0.025
r 60000_22000_M1 60000_24000_M1 0.025
r 60000_24000_M1 60000_26000_M1 0.025
r 60000_26000_M1 60000_28000_M1 0.025
r 60000_28000_M1 60000_30000_M1 0.025
r 60000_30000_M1 60000_32000_M1 0.025
r 60000_32000_M1 60000_34000_M1 0.025
r 60000_34000_M1 60000_36000_M1 0.025
r 60000_36000_M1 60000_38000_M1 0.025
r 60000_38000_M1 60000_40000_M1 0.025
r 60000_40000_M1 60000_42000_M1 0.025
r 60000_42000_M1 60000_44000_M1 0.025
r 60000_44000_M1 60000_46000_M1 0.025
r 60000_46000_M1 60000_48000_M1 0.025
r 60000_48000_M1 60000_50000_M1 0.025
r 60000_50000_M1 60000_52000_M1 0.025
r 60000_52000_M1 60000_54000_M1 0.025
r 60000_54000_M1 60000_56000_M1 0.025
r 60000_56000_M1 60000_58000_M1 0.025
r 60000_58000_M1 60000_60000_M1 0.025
r 60000_60000_M1 60000_62000_M1 0.025
r 60000_62000_M1 60000_64000_M1 0.025
r 60000_64000_M1 60000_66000_M1 0.025
r 60000_66000_M1 60000_68000_M1 0.025
r 60000_68000_M1 60000_70000_M1 0.025
r 60000_70000_M1 60000_72000_M1 0.025
r 60000_72000_M1 60000_74000_M1 0.025
r 60000_74000_M1 60000_76000_M1 0.025
r 60000_76000_M1 60000_78000_M1 0.025
r 60000_78000_M1 60000_80000_M1 0.025
r 60000_80000_M1 60000_82000_M1 0.025
r 60000_82000_M1 60000_84000_M1 0.025
r 60000_84000_M1 60000_86000_M1 0.025
r 60000_86000_M1 60000_88000_M1 0.025
r 60000_88000_M1 60000_90000_M1 0.025
r 60000_90000_M1 60000_92000_M1 0.025
r 60000_92000_M1 60000_94000_M1 0.025
r 60000_94000_M1 60000_96000_M1 0.025
r 60000_96000_M1 60000_98000_M1 0.025
r 60000_98000_M1 60000_100000_M1 0.025
r 62000_2000_M1 62000_4000_M1 0.025
r 62000_4000_M1 62000_6000_M1 0.025
r 62000_6000_M1 62000_8000_M1 0.025
r 62000_8000_M1 62000_10000_M1 0.025
r 62000_10000_M1 62000_12000_M1 0.025
r 62000_12000_M1 62000_14000_M1 0.025
r 62000_14000_M1 62000_16000_M1 0.025
r 62000_16000_M1 62000_18000_M1 0.025
r 62000_18000_M1 62000_20000_M1 0.025
r 62000_20000_M1 62000_22000_M1 0.025
r 62000_22000_M1 62000_24000_M1 0.025
r 62000_24000_M1 62000_26000_M1 0.025
r 62000_26000_M1 62000_28000_M1 0.025
r 62000_28000_M1 62000_30000_M1 0.025
r 62000_30000_M1 62000_32000_M1 0.025
r 62000_32000_M1 62000_34000_M1 0.025
r 62000_34000_M1 62000_36000_M1 0.025
r 62000_36000_M1 62000_38000_M1 0.025
r 62000_38000_M1 62000_40000_M1 0.025
r 62000_40000_M1 62000_42000_M1 0.025
r 62000_42000_M1 62000_44000_M1 0.025
r 62000_44000_M1 62000_46000_M1 0.025
r 62000_46000_M1 62000_48000_M1 0.025
r 62000_48000_M1 62000_50000_M1 0.025
r 62000_50000_M1 62000_52000_M1 0.025
r 62000_52000_M1 62000_54000_M1 0.025
r 62000_54000_M1 62000_56000_M1 0.025
r 62000_56000_M1 62000_58000_M1 0.025
r 62000_58000_M1 62000_60000_M1 0.025
r 62000_60000_M1 62000_62000_M1 0.025
r 62000_62000_M1 62000_64000_M1 0.025
r 62000_64000_M1 62000_66000_M1 0.025
r 62000_66000_M1 62000_68000_M1 0.025
r 62000_68000_M1 62000_70000_M1 0.025
r 62000_70000_M1 62000_72000_M1 0.025
r 62000_72000_M1 62000_74000_M1 0.025
r 62000_74000_M1 62000_76000_M1 0.025
r 62000_76000_M1 62000_78000_M1 0.025
r 62000_78000_M1 62000_80000_M1 0.025
r 62000_80000_M1 62000_82000_M1 0.025
r 62000_82000_M1 62000_84000_M1 0.025
r 62000_84000_M1 62000_86000_M1 0.025
r 62000_86000_M1 62000_88000_M1 0.025
r 62000_88000_M1 62000_90000_M1 0.025
r 62000_90000_M1 62000_92000_M1 0.025
r 62000_92000_M1 62000_94000_M1 0.025
r 62000_94000_M1 62000_96000_M1 0.025
r 62000_96000_M1 62000_98000_M1 0.025
r 62000_98000_M1 62000_100000_M1 0.025
r 64000_2000_M1 64000_4000_M1 0.025
r 64000_4000_M1 64000_6000_M1 0.025
r 64000_6000_M1 64000_8000_M1 0.025
r 64000_8000_M1 64000_10000_M1 0.025
r 64000_10000_M1 64000_12000_M1 0.025
r 64000_12000_M1 64000_14000_M1 0.025
r 64000_14000_M1 64000_16000_M1 0.025
r 64000_16000_M1 64000_18000_M1 0.025
r 64000_18000_M1 64000_20000_M1 0.025
r 64000_20000_M1 64000_22000_M1 0.025
r 64000_22000_M1 64000_24000_M1 0.025
r 64000_24000_M1 64000_26000_M1 0.025
r 64000_26000_M1 64000_28000_M1 0.025
r 64000_28000_M1 64000_30000_M1 0.025
r 64000_30000_M1 64000_32000_M1 0.025
r 64000_32000_M1 64000_34000_M1 0.025
r 64000_34000_M1 64000_36000_M1 0.025
r 64000_36000_M1 64000_38000_M1 0.025
r 64000_38000_M1 64000_40000_M1 0.025
r 64000_40000_M1 64000_42000_M1 0.025
r 64000_42000_M1 64000_44000_M1 0.025
r 64000_44000_M1 64000_46000_M1 0.025
r 64000_46000_M1 64000_48000_M1 0.025
r 64000_48000_M1 64000_50000_M1 0.025
r 64000_50000_M1 64000_52000_M1 0.025
r 64000_52000_M1 64000_54000_M1 0.025
r 64000_54000_M1 64000_56000_M1 0.025
r 64000_56000_M1 64000_58000_M1 0.025
r 64000_58000_M1 64000_60000_M1 0.025
r 64000_60000_M1 64000_62000_M1 0.025
r 64000_62000_M1 64000_64000_M1 0.025
r 64000_64000_M1 64000_66000_M1 0.025
r 64000_66000_M1 64000_68000_M1 0.025
r 64000_68000_M1 64000_70000_M1 0.025
r 64000_70000_M1 64000_72000_M1 0.025
r 64000_72000_M1 64000_74000_M1 0.025
r 64000_74000_M1 64000_76000_M1 0.025
r 64000_76000_M1 64000_78000_M1 0.025
r 64000_78000_M1 64000_80000_M1 0.025
r 64000_80000_M1 64000_82000_M1 0.025
r 64000_82000_M1 64000_84000_M1 0.025
r 64000_84000_M1 64000_86000_M1 0.025
r 64000_86000_M1 64000_88000_M1 0.025
r 64000_88000_M1 64000_90000_M1 0.025
r 64000_90000_M1 64000_92000_M1 0.025
r 64000_92000_M1 64000_94000_M1 0.025
r 64000_94000_M1 64000_96000_M1 0.025
r 64000_96000_M1 64000_98000_M1 0.025
r 64000_98000_M1 64000_100000_M1 0.025
r 66000_2000_M1 66000_4000_M1 0.025
r 66000_4000_M1 66000_6000_M1 0.025
r 66000_6000_M1 66000_8000_M1 0.025
r 66000_8000_M1 66000_10000_M1 0.025
r 66000_10000_M1 66000_12000_M1 0.025
r 66000_12000_M1 66000_14000_M1 0.025
r 66000_14000_M1 66000_16000_M1 0.025
r 66000_16000_M1 66000_18000_M1 0.025
r 66000_18000_M1 66000_20000_M1 0.025
r 66000_20000_M1 66000_22000_M1 0.025
r 66000_22000_M1 66000_24000_M1 0.025
r 66000_24000_M1 66000_26000_M1 0.025
r 66000_26000_M1 66000_28000_M1 0.025
r 66000_28000_M1 66000_30000_M1 0.025
r 66000_30000_M1 66000_32000_M1 0.025
r 66000_32000_M1 66000_34000_M1 0.025
r 66000_34000_M1 66000_36000_M1 0.025
r 66000_36000_M1 66000_38000_M1 0.025
r 66000_38000_M1 66000_40000_M1 0.025
r 66000_40000_M1 66000_42000_M1 0.025
r 66000_42000_M1 66000_44000_M1 0.025
r 66000_44000_M1 66000_46000_M1 0.025
r 66000_46000_M1 66000_48000_M1 0.025
r 66000_48000_M1 66000_50000_M1 0.025
r 66000_50000_M1 66000_52000_M1 0.025
r 66000_52000_M1 66000_54000_M1 0.025
r 66000_54000_M1 66000_56000_M1 0.025
r 66000_56000_M1 66000_58000_M1 0.025
r 66000_58000_M1 66000_60000_M1 0.025
r 66000_60000_M1 66000_62000_M1 0.025
r 66000_62000_M1 66000_64000_M1 0.025
r 66000_64000_M1 66000_66000_M1 0.025
r 66000_66000_M1 66000_68000_M1 0.025
r 66000_68000_M1 66000_70000_M1 0.025
r 66000_70000_M1 66000_72000_M1 0.025
r 66000_72000_M1 66000_74000_M1 0.025
r 66000_74000_M1 66000_76000_M1 0.025
r 66000_76000_M1 66000_78000_M1 0.025
r 66000_78000_M1 66000_80000_M1 0.025
r 66000_80000_M1 66000_82000_M1 0.025
r 66000_82000_M1 66000_84000_M1 0.025
r 66000_84000_M1 66000_86000_M1 0.025
r 66000_86000_M1 66000_88000_M1 0.025
r 66000_88000_M1 66000_90000_M1 0.025
r 66000_90000_M1 66000_92000_M1 0.025
r 66000_92000_M1 66000_94000_M1 0.025
r 66000_94000_M1 66000_96000_M1 0.025
r 66000_96000_M1 66000_98000_M1 0.025
r 66000_98000_M1 66000_100000_M1 0.025
r 68000_2000_M1 68000_4000_M1 0.025
r 68000_4000_M1 68000_6000_M1 0.025
r 68000_6000_M1 68000_8000_M1 0.025
r 68000_8000_M1 68000_10000_M1 0.025
r 68000_10000_M1 68000_12000_M1 0.025
r 68000_12000_M1 68000_14000_M1 0.025
r 68000_14000_M1 68000_16000_M1 0.025
r 68000_16000_M1 68000_18000_M1 0.025
r 68000_18000_M1 68000_20000_M1 0.025
r 68000_20000_M1 68000_22000_M1 0.025
r 68000_22000_M1 68000_24000_M1 0.025
r 68000_24000_M1 68000_26000_M1 0.025
r 68000_26000_M1 68000_28000_M1 0.025
r 68000_28000_M1 68000_30000_M1 0.025
r 68000_30000_M1 68000_32000_M1 0.025
r 68000_32000_M1 68000_34000_M1 0.025
r 68000_34000_M1 68000_36000_M1 0.025
r 68000_36000_M1 68000_38000_M1 0.025
r 68000_38000_M1 68000_40000_M1 0.025
r 68000_40000_M1 68000_42000_M1 0.025
r 68000_42000_M1 68000_44000_M1 0.025
r 68000_44000_M1 68000_46000_M1 0.025
r 68000_46000_M1 68000_48000_M1 0.025
r 68000_48000_M1 68000_50000_M1 0.025
r 68000_50000_M1 68000_52000_M1 0.025
r 68000_52000_M1 68000_54000_M1 0.025
r 68000_54000_M1 68000_56000_M1 0.025
r 68000_56000_M1 68000_58000_M1 0.025
r 68000_58000_M1 68000_60000_M1 0.025
r 68000_60000_M1 68000_62000_M1 0.025
r 68000_62000_M1 68000_64000_M1 0.025
r 68000_64000_M1 68000_66000_M1 0.025
r 68000_66000_M1 68000_68000_M1 0.025
r 68000_68000_M1 68000_70000_M1 0.025
r 68000_70000_M1 68000_72000_M1 0.025
r 68000_72000_M1 68000_74000_M1 0.025
r 68000_74000_M1 68000_76000_M1 0.025
r 68000_76000_M1 68000_78000_M1 0.025
r 68000_78000_M1 68000_80000_M1 0.025
r 68000_80000_M1 68000_82000_M1 0.025
r 68000_82000_M1 68000_84000_M1 0.025
r 68000_84000_M1 68000_86000_M1 0.025
r 68000_86000_M1 68000_88000_M1 0.025
r 68000_88000_M1 68000_90000_M1 0.025
r 68000_90000_M1 68000_92000_M1 0.025
r 68000_92000_M1 68000_94000_M1 0.025
r 68000_94000_M1 68000_96000_M1 0.025
r 68000_96000_M1 68000_98000_M1 0.025
r 68000_98000_M1 68000_100000_M1 0.025
r 70000_2000_M1 70000_4000_M1 0.025
r 70000_4000_M1 70000_6000_M1 0.025
r 70000_6000_M1 70000_8000_M1 0.025
r 70000_8000_M1 70000_10000_M1 0.025
r 70000_10000_M1 70000_12000_M1 0.025
r 70000_12000_M1 70000_14000_M1 0.025
r 70000_14000_M1 70000_16000_M1 0.025
r 70000_16000_M1 70000_18000_M1 0.025
r 70000_18000_M1 70000_20000_M1 0.025
r 70000_20000_M1 70000_22000_M1 0.025
r 70000_22000_M1 70000_24000_M1 0.025
r 70000_24000_M1 70000_26000_M1 0.025
r 70000_26000_M1 70000_28000_M1 0.025
r 70000_28000_M1 70000_30000_M1 0.025
r 70000_30000_M1 70000_32000_M1 0.025
r 70000_32000_M1 70000_34000_M1 0.025
r 70000_34000_M1 70000_36000_M1 0.025
r 70000_36000_M1 70000_38000_M1 0.025
r 70000_38000_M1 70000_40000_M1 0.025
r 70000_40000_M1 70000_42000_M1 0.025
r 70000_42000_M1 70000_44000_M1 0.025
r 70000_44000_M1 70000_46000_M1 0.025
r 70000_46000_M1 70000_48000_M1 0.025
r 70000_48000_M1 70000_50000_M1 0.025
r 70000_50000_M1 70000_52000_M1 0.025
r 70000_52000_M1 70000_54000_M1 0.025
r 70000_54000_M1 70000_56000_M1 0.025
r 70000_56000_M1 70000_58000_M1 0.025
r 70000_58000_M1 70000_60000_M1 0.025
r 70000_60000_M1 70000_62000_M1 0.025
r 70000_62000_M1 70000_64000_M1 0.025
r 70000_64000_M1 70000_66000_M1 0.025
r 70000_66000_M1 70000_68000_M1 0.025
r 70000_68000_M1 70000_70000_M1 0.025
r 70000_70000_M1 70000_72000_M1 0.025
r 70000_72000_M1 70000_74000_M1 0.025
r 70000_74000_M1 70000_76000_M1 0.025
r 70000_76000_M1 70000_78000_M1 0.025
r 70000_78000_M1 70000_80000_M1 0.025
r 70000_80000_M1 70000_82000_M1 0.025
r 70000_82000_M1 70000_84000_M1 0.025
r 70000_84000_M1 70000_86000_M1 0.025
r 70000_86000_M1 70000_88000_M1 0.025
r 70000_88000_M1 70000_90000_M1 0.025
r 70000_90000_M1 70000_92000_M1 0.025
r 70000_92000_M1 70000_94000_M1 0.025
r 70000_94000_M1 70000_96000_M1 0.025
r 70000_96000_M1 70000_98000_M1 0.025
r 70000_98000_M1 70000_100000_M1 0.025
r 72000_2000_M1 72000_4000_M1 0.025
r 72000_4000_M1 72000_6000_M1 0.025
r 72000_6000_M1 72000_8000_M1 0.025
r 72000_8000_M1 72000_10000_M1 0.025
r 72000_10000_M1 72000_12000_M1 0.025
r 72000_12000_M1 72000_14000_M1 0.025
r 72000_14000_M1 72000_16000_M1 0.025
r 72000_16000_M1 72000_18000_M1 0.025
r 72000_18000_M1 72000_20000_M1 0.025
r 72000_20000_M1 72000_22000_M1 0.025
r 72000_22000_M1 72000_24000_M1 0.025
r 72000_24000_M1 72000_26000_M1 0.025
r 72000_26000_M1 72000_28000_M1 0.025
r 72000_28000_M1 72000_30000_M1 0.025
r 72000_30000_M1 72000_32000_M1 0.025
r 72000_32000_M1 72000_34000_M1 0.025
r 72000_34000_M1 72000_36000_M1 0.025
r 72000_36000_M1 72000_38000_M1 0.025
r 72000_38000_M1 72000_40000_M1 0.025
r 72000_40000_M1 72000_42000_M1 0.025
r 72000_42000_M1 72000_44000_M1 0.025
r 72000_44000_M1 72000_46000_M1 0.025
r 72000_46000_M1 72000_48000_M1 0.025
r 72000_48000_M1 72000_50000_M1 0.025
r 72000_50000_M1 72000_52000_M1 0.025
r 72000_52000_M1 72000_54000_M1 0.025
r 72000_54000_M1 72000_56000_M1 0.025
r 72000_56000_M1 72000_58000_M1 0.025
r 72000_58000_M1 72000_60000_M1 0.025
r 72000_60000_M1 72000_62000_M1 0.025
r 72000_62000_M1 72000_64000_M1 0.025
r 72000_64000_M1 72000_66000_M1 0.025
r 72000_66000_M1 72000_68000_M1 0.025
r 72000_68000_M1 72000_70000_M1 0.025
r 72000_70000_M1 72000_72000_M1 0.025
r 72000_72000_M1 72000_74000_M1 0.025
r 72000_74000_M1 72000_76000_M1 0.025
r 72000_76000_M1 72000_78000_M1 0.025
r 72000_78000_M1 72000_80000_M1 0.025
r 72000_80000_M1 72000_82000_M1 0.025
r 72000_82000_M1 72000_84000_M1 0.025
r 72000_84000_M1 72000_86000_M1 0.025
r 72000_86000_M1 72000_88000_M1 0.025
r 72000_88000_M1 72000_90000_M1 0.025
r 72000_90000_M1 72000_92000_M1 0.025
r 72000_92000_M1 72000_94000_M1 0.025
r 72000_94000_M1 72000_96000_M1 0.025
r 72000_96000_M1 72000_98000_M1 0.025
r 72000_98000_M1 72000_100000_M1 0.025
r 74000_2000_M1 74000_4000_M1 0.025
r 74000_4000_M1 74000_6000_M1 0.025
r 74000_6000_M1 74000_8000_M1 0.025
r 74000_8000_M1 74000_10000_M1 0.025
r 74000_10000_M1 74000_12000_M1 0.025
r 74000_12000_M1 74000_14000_M1 0.025
r 74000_14000_M1 74000_16000_M1 0.025
r 74000_16000_M1 74000_18000_M1 0.025
r 74000_18000_M1 74000_20000_M1 0.025
r 74000_20000_M1 74000_22000_M1 0.025
r 74000_22000_M1 74000_24000_M1 0.025
r 74000_24000_M1 74000_26000_M1 0.025
r 74000_26000_M1 74000_28000_M1 0.025
r 74000_28000_M1 74000_30000_M1 0.025
r 74000_30000_M1 74000_32000_M1 0.025
r 74000_32000_M1 74000_34000_M1 0.025
r 74000_34000_M1 74000_36000_M1 0.025
r 74000_36000_M1 74000_38000_M1 0.025
r 74000_38000_M1 74000_40000_M1 0.025
r 74000_40000_M1 74000_42000_M1 0.025
r 74000_42000_M1 74000_44000_M1 0.025
r 74000_44000_M1 74000_46000_M1 0.025
r 74000_46000_M1 74000_48000_M1 0.025
r 74000_48000_M1 74000_50000_M1 0.025
r 74000_50000_M1 74000_52000_M1 0.025
r 74000_52000_M1 74000_54000_M1 0.025
r 74000_54000_M1 74000_56000_M1 0.025
r 74000_56000_M1 74000_58000_M1 0.025
r 74000_58000_M1 74000_60000_M1 0.025
r 74000_60000_M1 74000_62000_M1 0.025
r 74000_62000_M1 74000_64000_M1 0.025
r 74000_64000_M1 74000_66000_M1 0.025
r 74000_66000_M1 74000_68000_M1 0.025
r 74000_68000_M1 74000_70000_M1 0.025
r 74000_70000_M1 74000_72000_M1 0.025
r 74000_72000_M1 74000_74000_M1 0.025
r 74000_74000_M1 74000_76000_M1 0.025
r 74000_76000_M1 74000_78000_M1 0.025
r 74000_78000_M1 74000_80000_M1 0.025
r 74000_80000_M1 74000_82000_M1 0.025
r 74000_82000_M1 74000_84000_M1 0.025
r 74000_84000_M1 74000_86000_M1 0.025
r 74000_86000_M1 74000_88000_M1 0.025
r 74000_88000_M1 74000_90000_M1 0.025
r 74000_90000_M1 74000_92000_M1 0.025
r 74000_92000_M1 74000_94000_M1 0.025
r 74000_94000_M1 74000_96000_M1 0.025
r 74000_96000_M1 74000_98000_M1 0.025
r 74000_98000_M1 74000_100000_M1 0.025
r 76000_2000_M1 76000_4000_M1 0.025
r 76000_4000_M1 76000_6000_M1 0.025
r 76000_6000_M1 76000_8000_M1 0.025
r 76000_8000_M1 76000_10000_M1 0.025
r 76000_10000_M1 76000_12000_M1 0.025
r 76000_12000_M1 76000_14000_M1 0.025
r 76000_14000_M1 76000_16000_M1 0.025
r 76000_16000_M1 76000_18000_M1 0.025
r 76000_18000_M1 76000_20000_M1 0.025
r 76000_20000_M1 76000_22000_M1 0.025
r 76000_22000_M1 76000_24000_M1 0.025
r 76000_24000_M1 76000_26000_M1 0.025
r 76000_26000_M1 76000_28000_M1 0.025
r 76000_28000_M1 76000_30000_M1 0.025
r 76000_30000_M1 76000_32000_M1 0.025
r 76000_32000_M1 76000_34000_M1 0.025
r 76000_34000_M1 76000_36000_M1 0.025
r 76000_36000_M1 76000_38000_M1 0.025
r 76000_38000_M1 76000_40000_M1 0.025
r 76000_40000_M1 76000_42000_M1 0.025
r 76000_42000_M1 76000_44000_M1 0.025
r 76000_44000_M1 76000_46000_M1 0.025
r 76000_46000_M1 76000_48000_M1 0.025
r 76000_48000_M1 76000_50000_M1 0.025
r 76000_50000_M1 76000_52000_M1 0.025
r 76000_52000_M1 76000_54000_M1 0.025
r 76000_54000_M1 76000_56000_M1 0.025
r 76000_56000_M1 76000_58000_M1 0.025
r 76000_58000_M1 76000_60000_M1 0.025
r 76000_60000_M1 76000_62000_M1 0.025
r 76000_62000_M1 76000_64000_M1 0.025
r 76000_64000_M1 76000_66000_M1 0.025
r 76000_66000_M1 76000_68000_M1 0.025
r 76000_68000_M1 76000_70000_M1 0.025
r 76000_70000_M1 76000_72000_M1 0.025
r 76000_72000_M1 76000_74000_M1 0.025
r 76000_74000_M1 76000_76000_M1 0.025
r 76000_76000_M1 76000_78000_M1 0.025
r 76000_78000_M1 76000_80000_M1 0.025
r 76000_80000_M1 76000_82000_M1 0.025
r 76000_82000_M1 76000_84000_M1 0.025
r 76000_84000_M1 76000_86000_M1 0.025
r 76000_86000_M1 76000_88000_M1 0.025
r 76000_88000_M1 76000_90000_M1 0.025
r 76000_90000_M1 76000_92000_M1 0.025
r 76000_92000_M1 76000_94000_M1 0.025
r 76000_94000_M1 76000_96000_M1 0.025
r 76000_96000_M1 76000_98000_M1 0.025
r 76000_98000_M1 76000_100000_M1 0.025
r 78000_2000_M1 78000_4000_M1 0.025
r 78000_4000_M1 78000_6000_M1 0.025
r 78000_6000_M1 78000_8000_M1 0.025
r 78000_8000_M1 78000_10000_M1 0.025
r 78000_10000_M1 78000_12000_M1 0.025
r 78000_12000_M1 78000_14000_M1 0.025
r 78000_14000_M1 78000_16000_M1 0.025
r 78000_16000_M1 78000_18000_M1 0.025
r 78000_18000_M1 78000_20000_M1 0.025
r 78000_20000_M1 78000_22000_M1 0.025
r 78000_22000_M1 78000_24000_M1 0.025
r 78000_24000_M1 78000_26000_M1 0.025
r 78000_26000_M1 78000_28000_M1 0.025
r 78000_28000_M1 78000_30000_M1 0.025
r 78000_30000_M1 78000_32000_M1 0.025
r 78000_32000_M1 78000_34000_M1 0.025
r 78000_34000_M1 78000_36000_M1 0.025
r 78000_36000_M1 78000_38000_M1 0.025
r 78000_38000_M1 78000_40000_M1 0.025
r 78000_40000_M1 78000_42000_M1 0.025
r 78000_42000_M1 78000_44000_M1 0.025
r 78000_44000_M1 78000_46000_M1 0.025
r 78000_46000_M1 78000_48000_M1 0.025
r 78000_48000_M1 78000_50000_M1 0.025
r 78000_50000_M1 78000_52000_M1 0.025
r 78000_52000_M1 78000_54000_M1 0.025
r 78000_54000_M1 78000_56000_M1 0.025
r 78000_56000_M1 78000_58000_M1 0.025
r 78000_58000_M1 78000_60000_M1 0.025
r 78000_60000_M1 78000_62000_M1 0.025
r 78000_62000_M1 78000_64000_M1 0.025
r 78000_64000_M1 78000_66000_M1 0.025
r 78000_66000_M1 78000_68000_M1 0.025
r 78000_68000_M1 78000_70000_M1 0.025
r 78000_70000_M1 78000_72000_M1 0.025
r 78000_72000_M1 78000_74000_M1 0.025
r 78000_74000_M1 78000_76000_M1 0.025
r 78000_76000_M1 78000_78000_M1 0.025
r 78000_78000_M1 78000_80000_M1 0.025
r 78000_80000_M1 78000_82000_M1 0.025
r 78000_82000_M1 78000_84000_M1 0.025
r 78000_84000_M1 78000_86000_M1 0.025
r 78000_86000_M1 78000_88000_M1 0.025
r 78000_88000_M1 78000_90000_M1 0.025
r 78000_90000_M1 78000_92000_M1 0.025
r 78000_92000_M1 78000_94000_M1 0.025
r 78000_94000_M1 78000_96000_M1 0.025
r 78000_96000_M1 78000_98000_M1 0.025
r 78000_98000_M1 78000_100000_M1 0.025
r 80000_2000_M1 80000_4000_M1 0.025
r 80000_4000_M1 80000_6000_M1 0.025
r 80000_6000_M1 80000_8000_M1 0.025
r 80000_8000_M1 80000_10000_M1 0.025
r 80000_10000_M1 80000_12000_M1 0.025
r 80000_12000_M1 80000_14000_M1 0.025
r 80000_14000_M1 80000_16000_M1 0.025
r 80000_16000_M1 80000_18000_M1 0.025
r 80000_18000_M1 80000_20000_M1 0.025
r 80000_20000_M1 80000_22000_M1 0.025
r 80000_22000_M1 80000_24000_M1 0.025
r 80000_24000_M1 80000_26000_M1 0.025
r 80000_26000_M1 80000_28000_M1 0.025
r 80000_28000_M1 80000_30000_M1 0.025
r 80000_30000_M1 80000_32000_M1 0.025
r 80000_32000_M1 80000_34000_M1 0.025
r 80000_34000_M1 80000_36000_M1 0.025
r 80000_36000_M1 80000_38000_M1 0.025
r 80000_38000_M1 80000_40000_M1 0.025
r 80000_40000_M1 80000_42000_M1 0.025
r 80000_42000_M1 80000_44000_M1 0.025
r 80000_44000_M1 80000_46000_M1 0.025
r 80000_46000_M1 80000_48000_M1 0.025
r 80000_48000_M1 80000_50000_M1 0.025
r 80000_50000_M1 80000_52000_M1 0.025
r 80000_52000_M1 80000_54000_M1 0.025
r 80000_54000_M1 80000_56000_M1 0.025
r 80000_56000_M1 80000_58000_M1 0.025
r 80000_58000_M1 80000_60000_M1 0.025
r 80000_60000_M1 80000_62000_M1 0.025
r 80000_62000_M1 80000_64000_M1 0.025
r 80000_64000_M1 80000_66000_M1 0.025
r 80000_66000_M1 80000_68000_M1 0.025
r 80000_68000_M1 80000_70000_M1 0.025
r 80000_70000_M1 80000_72000_M1 0.025
r 80000_72000_M1 80000_74000_M1 0.025
r 80000_74000_M1 80000_76000_M1 0.025
r 80000_76000_M1 80000_78000_M1 0.025
r 80000_78000_M1 80000_80000_M1 0.025
r 80000_80000_M1 80000_82000_M1 0.025
r 80000_82000_M1 80000_84000_M1 0.025
r 80000_84000_M1 80000_86000_M1 0.025
r 80000_86000_M1 80000_88000_M1 0.025
r 80000_88000_M1 80000_90000_M1 0.025
r 80000_90000_M1 80000_92000_M1 0.025
r 80000_92000_M1 80000_94000_M1 0.025
r 80000_94000_M1 80000_96000_M1 0.025
r 80000_96000_M1 80000_98000_M1 0.025
r 80000_98000_M1 80000_100000_M1 0.025
r 82000_2000_M1 82000_4000_M1 0.025
r 82000_4000_M1 82000_6000_M1 0.025
r 82000_6000_M1 82000_8000_M1 0.025
r 82000_8000_M1 82000_10000_M1 0.025
r 82000_10000_M1 82000_12000_M1 0.025
r 82000_12000_M1 82000_14000_M1 0.025
r 82000_14000_M1 82000_16000_M1 0.025
r 82000_16000_M1 82000_18000_M1 0.025
r 82000_18000_M1 82000_20000_M1 0.025
r 82000_20000_M1 82000_22000_M1 0.025
r 82000_22000_M1 82000_24000_M1 0.025
r 82000_24000_M1 82000_26000_M1 0.025
r 82000_26000_M1 82000_28000_M1 0.025
r 82000_28000_M1 82000_30000_M1 0.025
r 82000_30000_M1 82000_32000_M1 0.025
r 82000_32000_M1 82000_34000_M1 0.025
r 82000_34000_M1 82000_36000_M1 0.025
r 82000_36000_M1 82000_38000_M1 0.025
r 82000_38000_M1 82000_40000_M1 0.025
r 82000_40000_M1 82000_42000_M1 0.025
r 82000_42000_M1 82000_44000_M1 0.025
r 82000_44000_M1 82000_46000_M1 0.025
r 82000_46000_M1 82000_48000_M1 0.025
r 82000_48000_M1 82000_50000_M1 0.025
r 82000_50000_M1 82000_52000_M1 0.025
r 82000_52000_M1 82000_54000_M1 0.025
r 82000_54000_M1 82000_56000_M1 0.025
r 82000_56000_M1 82000_58000_M1 0.025
r 82000_58000_M1 82000_60000_M1 0.025
r 82000_60000_M1 82000_62000_M1 0.025
r 82000_62000_M1 82000_64000_M1 0.025
r 82000_64000_M1 82000_66000_M1 0.025
r 82000_66000_M1 82000_68000_M1 0.025
r 82000_68000_M1 82000_70000_M1 0.025
r 82000_70000_M1 82000_72000_M1 0.025
r 82000_72000_M1 82000_74000_M1 0.025
r 82000_74000_M1 82000_76000_M1 0.025
r 82000_76000_M1 82000_78000_M1 0.025
r 82000_78000_M1 82000_80000_M1 0.025
r 82000_80000_M1 82000_82000_M1 0.025
r 82000_82000_M1 82000_84000_M1 0.025
r 82000_84000_M1 82000_86000_M1 0.025
r 82000_86000_M1 82000_88000_M1 0.025
r 82000_88000_M1 82000_90000_M1 0.025
r 82000_90000_M1 82000_92000_M1 0.025
r 82000_92000_M1 82000_94000_M1 0.025
r 82000_94000_M1 82000_96000_M1 0.025
r 82000_96000_M1 82000_98000_M1 0.025
r 82000_98000_M1 82000_100000_M1 0.025
r 84000_2000_M1 84000_4000_M1 0.025
r 84000_4000_M1 84000_6000_M1 0.025
r 84000_6000_M1 84000_8000_M1 0.025
r 84000_8000_M1 84000_10000_M1 0.025
r 84000_10000_M1 84000_12000_M1 0.025
r 84000_12000_M1 84000_14000_M1 0.025
r 84000_14000_M1 84000_16000_M1 0.025
r 84000_16000_M1 84000_18000_M1 0.025
r 84000_18000_M1 84000_20000_M1 0.025
r 84000_20000_M1 84000_22000_M1 0.025
r 84000_22000_M1 84000_24000_M1 0.025
r 84000_24000_M1 84000_26000_M1 0.025
r 84000_26000_M1 84000_28000_M1 0.025
r 84000_28000_M1 84000_30000_M1 0.025
r 84000_30000_M1 84000_32000_M1 0.025
r 84000_32000_M1 84000_34000_M1 0.025
r 84000_34000_M1 84000_36000_M1 0.025
r 84000_36000_M1 84000_38000_M1 0.025
r 84000_38000_M1 84000_40000_M1 0.025
r 84000_40000_M1 84000_42000_M1 0.025
r 84000_42000_M1 84000_44000_M1 0.025
r 84000_44000_M1 84000_46000_M1 0.025
r 84000_46000_M1 84000_48000_M1 0.025
r 84000_48000_M1 84000_50000_M1 0.025
r 84000_50000_M1 84000_52000_M1 0.025
r 84000_52000_M1 84000_54000_M1 0.025
r 84000_54000_M1 84000_56000_M1 0.025
r 84000_56000_M1 84000_58000_M1 0.025
r 84000_58000_M1 84000_60000_M1 0.025
r 84000_60000_M1 84000_62000_M1 0.025
r 84000_62000_M1 84000_64000_M1 0.025
r 84000_64000_M1 84000_66000_M1 0.025
r 84000_66000_M1 84000_68000_M1 0.025
r 84000_68000_M1 84000_70000_M1 0.025
r 84000_70000_M1 84000_72000_M1 0.025
r 84000_72000_M1 84000_74000_M1 0.025
r 84000_74000_M1 84000_76000_M1 0.025
r 84000_76000_M1 84000_78000_M1 0.025
r 84000_78000_M1 84000_80000_M1 0.025
r 84000_80000_M1 84000_82000_M1 0.025
r 84000_82000_M1 84000_84000_M1 0.025
r 84000_84000_M1 84000_86000_M1 0.025
r 84000_86000_M1 84000_88000_M1 0.025
r 84000_88000_M1 84000_90000_M1 0.025
r 84000_90000_M1 84000_92000_M1 0.025
r 84000_92000_M1 84000_94000_M1 0.025
r 84000_94000_M1 84000_96000_M1 0.025
r 84000_96000_M1 84000_98000_M1 0.025
r 84000_98000_M1 84000_100000_M1 0.025
r 86000_2000_M1 86000_4000_M1 0.025
r 86000_4000_M1 86000_6000_M1 0.025
r 86000_6000_M1 86000_8000_M1 0.025
r 86000_8000_M1 86000_10000_M1 0.025
r 86000_10000_M1 86000_12000_M1 0.025
r 86000_12000_M1 86000_14000_M1 0.025
r 86000_14000_M1 86000_16000_M1 0.025
r 86000_16000_M1 86000_18000_M1 0.025
r 86000_18000_M1 86000_20000_M1 0.025
r 86000_20000_M1 86000_22000_M1 0.025
r 86000_22000_M1 86000_24000_M1 0.025
r 86000_24000_M1 86000_26000_M1 0.025
r 86000_26000_M1 86000_28000_M1 0.025
r 86000_28000_M1 86000_30000_M1 0.025
r 86000_30000_M1 86000_32000_M1 0.025
r 86000_32000_M1 86000_34000_M1 0.025
r 86000_34000_M1 86000_36000_M1 0.025
r 86000_36000_M1 86000_38000_M1 0.025
r 86000_38000_M1 86000_40000_M1 0.025
r 86000_40000_M1 86000_42000_M1 0.025
r 86000_42000_M1 86000_44000_M1 0.025
r 86000_44000_M1 86000_46000_M1 0.025
r 86000_46000_M1 86000_48000_M1 0.025
r 86000_48000_M1 86000_50000_M1 0.025
r 86000_50000_M1 86000_52000_M1 0.025
r 86000_52000_M1 86000_54000_M1 0.025
r 86000_54000_M1 86000_56000_M1 0.025
r 86000_56000_M1 86000_58000_M1 0.025
r 86000_58000_M1 86000_60000_M1 0.025
r 86000_60000_M1 86000_62000_M1 0.025
r 86000_62000_M1 86000_64000_M1 0.025
r 86000_64000_M1 86000_66000_M1 0.025
r 86000_66000_M1 86000_68000_M1 0.025
r 86000_68000_M1 86000_70000_M1 0.025
r 86000_70000_M1 86000_72000_M1 0.025
r 86000_72000_M1 86000_74000_M1 0.025
r 86000_74000_M1 86000_76000_M1 0.025
r 86000_76000_M1 86000_78000_M1 0.025
r 86000_78000_M1 86000_80000_M1 0.025
r 86000_80000_M1 86000_82000_M1 0.025
r 86000_82000_M1 86000_84000_M1 0.025
r 86000_84000_M1 86000_86000_M1 0.025
r 86000_86000_M1 86000_88000_M1 0.025
r 86000_88000_M1 86000_90000_M1 0.025
r 86000_90000_M1 86000_92000_M1 0.025
r 86000_92000_M1 86000_94000_M1 0.025
r 86000_94000_M1 86000_96000_M1 0.025
r 86000_96000_M1 86000_98000_M1 0.025
r 86000_98000_M1 86000_100000_M1 0.025
r 88000_2000_M1 88000_4000_M1 0.025
r 88000_4000_M1 88000_6000_M1 0.025
r 88000_6000_M1 88000_8000_M1 0.025
r 88000_8000_M1 88000_10000_M1 0.025
r 88000_10000_M1 88000_12000_M1 0.025
r 88000_12000_M1 88000_14000_M1 0.025
r 88000_14000_M1 88000_16000_M1 0.025
r 88000_16000_M1 88000_18000_M1 0.025
r 88000_18000_M1 88000_20000_M1 0.025
r 88000_20000_M1 88000_22000_M1 0.025
r 88000_22000_M1 88000_24000_M1 0.025
r 88000_24000_M1 88000_26000_M1 0.025
r 88000_26000_M1 88000_28000_M1 0.025
r 88000_28000_M1 88000_30000_M1 0.025
r 88000_30000_M1 88000_32000_M1 0.025
r 88000_32000_M1 88000_34000_M1 0.025
r 88000_34000_M1 88000_36000_M1 0.025
r 88000_36000_M1 88000_38000_M1 0.025
r 88000_38000_M1 88000_40000_M1 0.025
r 88000_40000_M1 88000_42000_M1 0.025
r 88000_42000_M1 88000_44000_M1 0.025
r 88000_44000_M1 88000_46000_M1 0.025
r 88000_46000_M1 88000_48000_M1 0.025
r 88000_48000_M1 88000_50000_M1 0.025
r 88000_50000_M1 88000_52000_M1 0.025
r 88000_52000_M1 88000_54000_M1 0.025
r 88000_54000_M1 88000_56000_M1 0.025
r 88000_56000_M1 88000_58000_M1 0.025
r 88000_58000_M1 88000_60000_M1 0.025
r 88000_60000_M1 88000_62000_M1 0.025
r 88000_62000_M1 88000_64000_M1 0.025
r 88000_64000_M1 88000_66000_M1 0.025
r 88000_66000_M1 88000_68000_M1 0.025
r 88000_68000_M1 88000_70000_M1 0.025
r 88000_70000_M1 88000_72000_M1 0.025
r 88000_72000_M1 88000_74000_M1 0.025
r 88000_74000_M1 88000_76000_M1 0.025
r 88000_76000_M1 88000_78000_M1 0.025
r 88000_78000_M1 88000_80000_M1 0.025
r 88000_80000_M1 88000_82000_M1 0.025
r 88000_82000_M1 88000_84000_M1 0.025
r 88000_84000_M1 88000_86000_M1 0.025
r 88000_86000_M1 88000_88000_M1 0.025
r 88000_88000_M1 88000_90000_M1 0.025
r 88000_90000_M1 88000_92000_M1 0.025
r 88000_92000_M1 88000_94000_M1 0.025
r 88000_94000_M1 88000_96000_M1 0.025
r 88000_96000_M1 88000_98000_M1 0.025
r 88000_98000_M1 88000_100000_M1 0.025
r 90000_2000_M1 90000_4000_M1 0.025
r 90000_4000_M1 90000_6000_M1 0.025
r 90000_6000_M1 90000_8000_M1 0.025
r 90000_8000_M1 90000_10000_M1 0.025
r 90000_10000_M1 90000_12000_M1 0.025
r 90000_12000_M1 90000_14000_M1 0.025
r 90000_14000_M1 90000_16000_M1 0.025
r 90000_16000_M1 90000_18000_M1 0.025
r 90000_18000_M1 90000_20000_M1 0.025
r 90000_20000_M1 90000_22000_M1 0.025
r 90000_22000_M1 90000_24000_M1 0.025
r 90000_24000_M1 90000_26000_M1 0.025
r 90000_26000_M1 90000_28000_M1 0.025
r 90000_28000_M1 90000_30000_M1 0.025
r 90000_30000_M1 90000_32000_M1 0.025
r 90000_32000_M1 90000_34000_M1 0.025
r 90000_34000_M1 90000_36000_M1 0.025
r 90000_36000_M1 90000_38000_M1 0.025
r 90000_38000_M1 90000_40000_M1 0.025
r 90000_40000_M1 90000_42000_M1 0.025
r 90000_42000_M1 90000_44000_M1 0.025
r 90000_44000_M1 90000_46000_M1 0.025
r 90000_46000_M1 90000_48000_M1 0.025
r 90000_48000_M1 90000_50000_M1 0.025
r 90000_50000_M1 90000_52000_M1 0.025
r 90000_52000_M1 90000_54000_M1 0.025
r 90000_54000_M1 90000_56000_M1 0.025
r 90000_56000_M1 90000_58000_M1 0.025
r 90000_58000_M1 90000_60000_M1 0.025
r 90000_60000_M1 90000_62000_M1 0.025
r 90000_62000_M1 90000_64000_M1 0.025
r 90000_64000_M1 90000_66000_M1 0.025
r 90000_66000_M1 90000_68000_M1 0.025
r 90000_68000_M1 90000_70000_M1 0.025
r 90000_70000_M1 90000_72000_M1 0.025
r 90000_72000_M1 90000_74000_M1 0.025
r 90000_74000_M1 90000_76000_M1 0.025
r 90000_76000_M1 90000_78000_M1 0.025
r 90000_78000_M1 90000_80000_M1 0.025
r 90000_80000_M1 90000_82000_M1 0.025
r 90000_82000_M1 90000_84000_M1 0.025
r 90000_84000_M1 90000_86000_M1 0.025
r 90000_86000_M1 90000_88000_M1 0.025
r 90000_88000_M1 90000_90000_M1 0.025
r 90000_90000_M1 90000_92000_M1 0.025
r 90000_92000_M1 90000_94000_M1 0.025
r 90000_94000_M1 90000_96000_M1 0.025
r 90000_96000_M1 90000_98000_M1 0.025
r 90000_98000_M1 90000_100000_M1 0.025
r 92000_2000_M1 92000_4000_M1 0.025
r 92000_4000_M1 92000_6000_M1 0.025
r 92000_6000_M1 92000_8000_M1 0.025
r 92000_8000_M1 92000_10000_M1 0.025
r 92000_10000_M1 92000_12000_M1 0.025
r 92000_12000_M1 92000_14000_M1 0.025
r 92000_14000_M1 92000_16000_M1 0.025
r 92000_16000_M1 92000_18000_M1 0.025
r 92000_18000_M1 92000_20000_M1 0.025
r 92000_20000_M1 92000_22000_M1 0.025
r 92000_22000_M1 92000_24000_M1 0.025
r 92000_24000_M1 92000_26000_M1 0.025
r 92000_26000_M1 92000_28000_M1 0.025
r 92000_28000_M1 92000_30000_M1 0.025
r 92000_30000_M1 92000_32000_M1 0.025
r 92000_32000_M1 92000_34000_M1 0.025
r 92000_34000_M1 92000_36000_M1 0.025
r 92000_36000_M1 92000_38000_M1 0.025
r 92000_38000_M1 92000_40000_M1 0.025
r 92000_40000_M1 92000_42000_M1 0.025
r 92000_42000_M1 92000_44000_M1 0.025
r 92000_44000_M1 92000_46000_M1 0.025
r 92000_46000_M1 92000_48000_M1 0.025
r 92000_48000_M1 92000_50000_M1 0.025
r 92000_50000_M1 92000_52000_M1 0.025
r 92000_52000_M1 92000_54000_M1 0.025
r 92000_54000_M1 92000_56000_M1 0.025
r 92000_56000_M1 92000_58000_M1 0.025
r 92000_58000_M1 92000_60000_M1 0.025
r 92000_60000_M1 92000_62000_M1 0.025
r 92000_62000_M1 92000_64000_M1 0.025
r 92000_64000_M1 92000_66000_M1 0.025
r 92000_66000_M1 92000_68000_M1 0.025
r 92000_68000_M1 92000_70000_M1 0.025
r 92000_70000_M1 92000_72000_M1 0.025
r 92000_72000_M1 92000_74000_M1 0.025
r 92000_74000_M1 92000_76000_M1 0.025
r 92000_76000_M1 92000_78000_M1 0.025
r 92000_78000_M1 92000_80000_M1 0.025
r 92000_80000_M1 92000_82000_M1 0.025
r 92000_82000_M1 92000_84000_M1 0.025
r 92000_84000_M1 92000_86000_M1 0.025
r 92000_86000_M1 92000_88000_M1 0.025
r 92000_88000_M1 92000_90000_M1 0.025
r 92000_90000_M1 92000_92000_M1 0.025
r 92000_92000_M1 92000_94000_M1 0.025
r 92000_94000_M1 92000_96000_M1 0.025
r 92000_96000_M1 92000_98000_M1 0.025
r 92000_98000_M1 92000_100000_M1 0.025
r 94000_2000_M1 94000_4000_M1 0.025
r 94000_4000_M1 94000_6000_M1 0.025
r 94000_6000_M1 94000_8000_M1 0.025
r 94000_8000_M1 94000_10000_M1 0.025
r 94000_10000_M1 94000_12000_M1 0.025
r 94000_12000_M1 94000_14000_M1 0.025
r 94000_14000_M1 94000_16000_M1 0.025
r 94000_16000_M1 94000_18000_M1 0.025
r 94000_18000_M1 94000_20000_M1 0.025
r 94000_20000_M1 94000_22000_M1 0.025
r 94000_22000_M1 94000_24000_M1 0.025
r 94000_24000_M1 94000_26000_M1 0.025
r 94000_26000_M1 94000_28000_M1 0.025
r 94000_28000_M1 94000_30000_M1 0.025
r 94000_30000_M1 94000_32000_M1 0.025
r 94000_32000_M1 94000_34000_M1 0.025
r 94000_34000_M1 94000_36000_M1 0.025
r 94000_36000_M1 94000_38000_M1 0.025
r 94000_38000_M1 94000_40000_M1 0.025
r 94000_40000_M1 94000_42000_M1 0.025
r 94000_42000_M1 94000_44000_M1 0.025
r 94000_44000_M1 94000_46000_M1 0.025
r 94000_46000_M1 94000_48000_M1 0.025
r 94000_48000_M1 94000_50000_M1 0.025
r 94000_50000_M1 94000_52000_M1 0.025
r 94000_52000_M1 94000_54000_M1 0.025
r 94000_54000_M1 94000_56000_M1 0.025
r 94000_56000_M1 94000_58000_M1 0.025
r 94000_58000_M1 94000_60000_M1 0.025
r 94000_60000_M1 94000_62000_M1 0.025
r 94000_62000_M1 94000_64000_M1 0.025
r 94000_64000_M1 94000_66000_M1 0.025
r 94000_66000_M1 94000_68000_M1 0.025
r 94000_68000_M1 94000_70000_M1 0.025
r 94000_70000_M1 94000_72000_M1 0.025
r 94000_72000_M1 94000_74000_M1 0.025
r 94000_74000_M1 94000_76000_M1 0.025
r 94000_76000_M1 94000_78000_M1 0.025
r 94000_78000_M1 94000_80000_M1 0.025
r 94000_80000_M1 94000_82000_M1 0.025
r 94000_82000_M1 94000_84000_M1 0.025
r 94000_84000_M1 94000_86000_M1 0.025
r 94000_86000_M1 94000_88000_M1 0.025
r 94000_88000_M1 94000_90000_M1 0.025
r 94000_90000_M1 94000_92000_M1 0.025
r 94000_92000_M1 94000_94000_M1 0.025
r 94000_94000_M1 94000_96000_M1 0.025
r 94000_96000_M1 94000_98000_M1 0.025
r 94000_98000_M1 94000_100000_M1 0.025
r 96000_2000_M1 96000_4000_M1 0.025
r 96000_4000_M1 96000_6000_M1 0.025
r 96000_6000_M1 96000_8000_M1 0.025
r 96000_8000_M1 96000_10000_M1 0.025
r 96000_10000_M1 96000_12000_M1 0.025
r 96000_12000_M1 96000_14000_M1 0.025
r 96000_14000_M1 96000_16000_M1 0.025
r 96000_16000_M1 96000_18000_M1 0.025
r 96000_18000_M1 96000_20000_M1 0.025
r 96000_20000_M1 96000_22000_M1 0.025
r 96000_22000_M1 96000_24000_M1 0.025
r 96000_24000_M1 96000_26000_M1 0.025
r 96000_26000_M1 96000_28000_M1 0.025
r 96000_28000_M1 96000_30000_M1 0.025
r 96000_30000_M1 96000_32000_M1 0.025
r 96000_32000_M1 96000_34000_M1 0.025
r 96000_34000_M1 96000_36000_M1 0.025
r 96000_36000_M1 96000_38000_M1 0.025
r 96000_38000_M1 96000_40000_M1 0.025
r 96000_40000_M1 96000_42000_M1 0.025
r 96000_42000_M1 96000_44000_M1 0.025
r 96000_44000_M1 96000_46000_M1 0.025
r 96000_46000_M1 96000_48000_M1 0.025
r 96000_48000_M1 96000_50000_M1 0.025
r 96000_50000_M1 96000_52000_M1 0.025
r 96000_52000_M1 96000_54000_M1 0.025
r 96000_54000_M1 96000_56000_M1 0.025
r 96000_56000_M1 96000_58000_M1 0.025
r 96000_58000_M1 96000_60000_M1 0.025
r 96000_60000_M1 96000_62000_M1 0.025
r 96000_62000_M1 96000_64000_M1 0.025
r 96000_64000_M1 96000_66000_M1 0.025
r 96000_66000_M1 96000_68000_M1 0.025
r 96000_68000_M1 96000_70000_M1 0.025
r 96000_70000_M1 96000_72000_M1 0.025
r 96000_72000_M1 96000_74000_M1 0.025
r 96000_74000_M1 96000_76000_M1 0.025
r 96000_76000_M1 96000_78000_M1 0.025
r 96000_78000_M1 96000_80000_M1 0.025
r 96000_80000_M1 96000_82000_M1 0.025
r 96000_82000_M1 96000_84000_M1 0.025
r 96000_84000_M1 96000_86000_M1 0.025
r 96000_86000_M1 96000_88000_M1 0.025
r 96000_88000_M1 96000_90000_M1 0.025
r 96000_90000_M1 96000_92000_M1 0.025
r 96000_92000_M1 96000_94000_M1 0.025
r 96000_94000_M1 96000_96000_M1 0.025
r 96000_96000_M1 96000_98000_M1 0.025
r 96000_98000_M1 96000_100000_M1 0.025
r 98000_2000_M1 98000_4000_M1 0.025
r 98000_4000_M1 98000_6000_M1 0.025
r 98000_6000_M1 98000_8000_M1 0.025
r 98000_8000_M1 98000_10000_M1 0.025
r 98000_10000_M1 98000_12000_M1 0.025
r 98000_12000_M1 98000_14000_M1 0.025
r 98000_14000_M1 98000_16000_M1 0.025
r 98000_16000_M1 98000_18000_M1 0.025
r 98000_18000_M1 98000_20000_M1 0.025
r 98000_20000_M1 98000_22000_M1 0.025
r 98000_22000_M1 98000_24000_M1 0.025
r 98000_24000_M1 98000_26000_M1 0.025
r 98000_26000_M1 98000_28000_M1 0.025
r 98000_28000_M1 98000_30000_M1 0.025
r 98000_30000_M1 98000_32000_M1 0.025
r 98000_32000_M1 98000_34000_M1 0.025
r 98000_34000_M1 98000_36000_M1 0.025
r 98000_36000_M1 98000_38000_M1 0.025
r 98000_38000_M1 98000_40000_M1 0.025
r 98000_40000_M1 98000_42000_M1 0.025
r 98000_42000_M1 98000_44000_M1 0.025
r 98000_44000_M1 98000_46000_M1 0.025
r 98000_46000_M1 98000_48000_M1 0.025
r 98000_48000_M1 98000_50000_M1 0.025
r 98000_50000_M1 98000_52000_M1 0.025
r 98000_52000_M1 98000_54000_M1 0.025
r 98000_54000_M1 98000_56000_M1 0.025
r 98000_56000_M1 98000_58000_M1 0.025
r 98000_58000_M1 98000_60000_M1 0.025
r 98000_60000_M1 98000_62000_M1 0.025
r 98000_62000_M1 98000_64000_M1 0.025
r 98000_64000_M1 98000_66000_M1 0.025
r 98000_66000_M1 98000_68000_M1 0.025
r 98000_68000_M1 98000_70000_M1 0.025
r 98000_70000_M1 98000_72000_M1 0.025
r 98000_72000_M1 98000_74000_M1 0.025
r 98000_74000_M1 98000_76000_M1 0.025
r 98000_76000_M1 98000_78000_M1 0.025
r 98000_78000_M1 98000_80000_M1 0.025
r 98000_80000_M1 98000_82000_M1 0.025
r 98000_82000_M1 98000_84000_M1 0.025
r 98000_84000_M1 98000_86000_M1 0.025
r 98000_86000_M1 98000_88000_M1 0.025
r 98000_88000_M1 98000_90000_M1 0.025
r 98000_90000_M1 98000_92000_M1 0.025
r 98000_92000_M1 98000_94000_M1 0.025
r 98000_94000_M1 98000_96000_M1 0.025
r 98000_96000_M1 98000_98000_M1 0.025
r 98000_98000_M1 98000_100000_M1 0.025
r 100000_2000_M1 100000_4000_M1 0.025
r 100000_4000_M1 100000_6000_M1 0.025
r 100000_6000_M1 100000_8000_M1 0.025
r 100000_8000_M1 100000_10000_M1 0.025
r 100000_10000_M1 100000_12000_M1 0.025
r 100000_12000_M1 100000_14000_M1 0.025
r 100000_14000_M1 100000_16000_M1 0.025
r 100000_16000_M1 100000_18000_M1 0.025
r 100000_18000_M1 100000_20000_M1 0.025
r 100000_20000_M1 100000_22000_M1 0.025
r 100000_22000_M1 100000_24000_M1 0.025
r 100000_24000_M1 100000_26000_M1 0.025
r 100000_26000_M1 100000_28000_M1 0.025
r 100000_28000_M1 100000_30000_M1 0.025
r 100000_30000_M1 100000_32000_M1 0.025
r 100000_32000_M1 100000_34000_M1 0.025
r 100000_34000_M1 100000_36000_M1 0.025
r 100000_36000_M1 100000_38000_M1 0.025
r 100000_38000_M1 100000_40000_M1 0.025
r 100000_40000_M1 100000_42000_M1 0.025
r 100000_42000_M1 100000_44000_M1 0.025
r 100000_44000_M1 100000_46000_M1 0.025
r 100000_46000_M1 100000_48000_M1 0.025
r 100000_48000_M1 100000_50000_M1 0.025
r 100000_50000_M1 100000_52000_M1 0.025
r 100000_52000_M1 100000_54000_M1 0.025
r 100000_54000_M1 100000_56000_M1 0.025
r 100000_56000_M1 100000_58000_M1 0.025
r 100000_58000_M1 100000_60000_M1 0.025
r 100000_60000_M1 100000_62000_M1 0.025
r 100000_62000_M1 100000_64000_M1 0.025
r 100000_64000_M1 100000_66000_M1 0.025
r 100000_66000_M1 100000_68000_M1 0.025
r 100000_68000_M1 100000_70000_M1 0.025
r 100000_70000_M1 100000_72000_M1 0.025
r 100000_72000_M1 100000_74000_M1 0.025
r 100000_74000_M1 100000_76000_M1 0.025
r 100000_76000_M1 100000_78000_M1 0.025
r 100000_78000_M1 100000_80000_M1 0.025
r 100000_80000_M1 100000_82000_M1 0.025
r 100000_82000_M1 100000_84000_M1 0.025
r 100000_84000_M1 100000_86000_M1 0.025
r 100000_86000_M1 100000_88000_M1 0.025
r 100000_88000_M1 100000_90000_M1 0.025
r 100000_90000_M1 100000_92000_M1 0.025
r 100000_92000_M1 100000_94000_M1 0.025
r 100000_94000_M1 100000_96000_M1 0.025
r 100000_96000_M1 100000_98000_M1 0.025
r 100000_98000_M1 100000_100000_M1 0.025

* ============================================================================
* Layer M2 - 50x50 grid
* ============================================================================

* M2 Horizontal resistors
r 2000_2000_M2 4000_2000_M2 0.018
r 4000_2000_M2 6000_2000_M2 0.018
r 6000_2000_M2 8000_2000_M2 0.018
r 8000_2000_M2 10000_2000_M2 0.018
r 10000_2000_M2 12000_2000_M2 0.018
r 12000_2000_M2 14000_2000_M2 0.018
r 14000_2000_M2 16000_2000_M2 0.018
r 16000_2000_M2 18000_2000_M2 0.018
r 18000_2000_M2 20000_2000_M2 0.018
r 20000_2000_M2 22000_2000_M2 0.018
r 22000_2000_M2 24000_2000_M2 0.018
r 24000_2000_M2 26000_2000_M2 0.018
r 26000_2000_M2 28000_2000_M2 0.018
r 28000_2000_M2 30000_2000_M2 0.018
r 30000_2000_M2 32000_2000_M2 0.018
r 32000_2000_M2 34000_2000_M2 0.018
r 34000_2000_M2 36000_2000_M2 0.018
r 36000_2000_M2 38000_2000_M2 0.018
r 38000_2000_M2 40000_2000_M2 0.018
r 40000_2000_M2 42000_2000_M2 0.018
r 42000_2000_M2 44000_2000_M2 0.018
r 44000_2000_M2 46000_2000_M2 0.018
r 46000_2000_M2 48000_2000_M2 0.018
r 48000_2000_M2 50000_2000_M2 0.018
r 50000_2000_M2 52000_2000_M2 0.018
r 52000_2000_M2 54000_2000_M2 0.018
r 54000_2000_M2 56000_2000_M2 0.018
r 56000_2000_M2 58000_2000_M2 0.018
r 58000_2000_M2 60000_2000_M2 0.018
r 60000_2000_M2 62000_2000_M2 0.018
r 62000_2000_M2 64000_2000_M2 0.018
r 64000_2000_M2 66000_2000_M2 0.018
r 66000_2000_M2 68000_2000_M2 0.018
r 68000_2000_M2 70000_2000_M2 0.018
r 70000_2000_M2 72000_2000_M2 0.018
r 72000_2000_M2 74000_2000_M2 0.018
r 74000_2000_M2 76000_2000_M2 0.018
r 76000_2000_M2 78000_2000_M2 0.018
r 78000_2000_M2 80000_2000_M2 0.018
r 80000_2000_M2 82000_2000_M2 0.018
r 82000_2000_M2 84000_2000_M2 0.018
r 84000_2000_M2 86000_2000_M2 0.018
r 86000_2000_M2 88000_2000_M2 0.018
r 88000_2000_M2 90000_2000_M2 0.018
r 90000_2000_M2 92000_2000_M2 0.018
r 92000_2000_M2 94000_2000_M2 0.018
r 94000_2000_M2 96000_2000_M2 0.018
r 96000_2000_M2 98000_2000_M2 0.018
r 98000_2000_M2 100000_2000_M2 0.018
r 2000_4000_M2 4000_4000_M2 0.018
r 4000_4000_M2 6000_4000_M2 0.018
r 6000_4000_M2 8000_4000_M2 0.018
r 8000_4000_M2 10000_4000_M2 0.018
r 10000_4000_M2 12000_4000_M2 0.018
r 12000_4000_M2 14000_4000_M2 0.018
r 14000_4000_M2 16000_4000_M2 0.018
r 16000_4000_M2 18000_4000_M2 0.018
r 18000_4000_M2 20000_4000_M2 0.018
r 20000_4000_M2 22000_4000_M2 0.018
r 22000_4000_M2 24000_4000_M2 0.018
r 24000_4000_M2 26000_4000_M2 0.018
r 26000_4000_M2 28000_4000_M2 0.018
r 28000_4000_M2 30000_4000_M2 0.018
r 30000_4000_M2 32000_4000_M2 0.018
r 32000_4000_M2 34000_4000_M2 0.018
r 34000_4000_M2 36000_4000_M2 0.018
r 36000_4000_M2 38000_4000_M2 0.018
r 38000_4000_M2 40000_4000_M2 0.018
r 40000_4000_M2 42000_4000_M2 0.018
r 42000_4000_M2 44000_4000_M2 0.018
r 44000_4000_M2 46000_4000_M2 0.018
r 46000_4000_M2 48000_4000_M2 0.018
r 48000_4000_M2 50000_4000_M2 0.018
r 50000_4000_M2 52000_4000_M2 0.018
r 52000_4000_M2 54000_4000_M2 0.018
r 54000_4000_M2 56000_4000_M2 0.018
r 56000_4000_M2 58000_4000_M2 0.018
r 58000_4000_M2 60000_4000_M2 0.018
r 60000_4000_M2 62000_4000_M2 0.018
r 62000_4000_M2 64000_4000_M2 0.018
r 64000_4000_M2 66000_4000_M2 0.018
r 66000_4000_M2 68000_4000_M2 0.018
r 68000_4000_M2 70000_4000_M2 0.018
r 70000_4000_M2 72000_4000_M2 0.018
r 72000_4000_M2 74000_4000_M2 0.018
r 74000_4000_M2 76000_4000_M2 0.018
r 76000_4000_M2 78000_4000_M2 0.018
r 78000_4000_M2 80000_4000_M2 0.018
r 80000_4000_M2 82000_4000_M2 0.018
r 82000_4000_M2 84000_4000_M2 0.018
r 84000_4000_M2 86000_4000_M2 0.018
r 86000_4000_M2 88000_4000_M2 0.018
r 88000_4000_M2 90000_4000_M2 0.018
r 90000_4000_M2 92000_4000_M2 0.018
r 92000_4000_M2 94000_4000_M2 0.018
r 94000_4000_M2 96000_4000_M2 0.018
r 96000_4000_M2 98000_4000_M2 0.018
r 98000_4000_M2 100000_4000_M2 0.018
r 2000_6000_M2 4000_6000_M2 0.018
r 4000_6000_M2 6000_6000_M2 0.018
r 6000_6000_M2 8000_6000_M2 0.018
r 8000_6000_M2 10000_6000_M2 0.018
r 10000_6000_M2 12000_6000_M2 0.018
r 12000_6000_M2 14000_6000_M2 0.018
r 14000_6000_M2 16000_6000_M2 0.018
r 16000_6000_M2 18000_6000_M2 0.018
r 18000_6000_M2 20000_6000_M2 0.018
r 20000_6000_M2 22000_6000_M2 0.018
r 22000_6000_M2 24000_6000_M2 0.018
r 24000_6000_M2 26000_6000_M2 0.018
r 26000_6000_M2 28000_6000_M2 0.018
r 28000_6000_M2 30000_6000_M2 0.018
r 30000_6000_M2 32000_6000_M2 0.018
r 32000_6000_M2 34000_6000_M2 0.018
r 34000_6000_M2 36000_6000_M2 0.018
r 36000_6000_M2 38000_6000_M2 0.018
r 38000_6000_M2 40000_6000_M2 0.018
r 40000_6000_M2 42000_6000_M2 0.018
r 42000_6000_M2 44000_6000_M2 0.018
r 44000_6000_M2 46000_6000_M2 0.018
r 46000_6000_M2 48000_6000_M2 0.018
r 48000_6000_M2 50000_6000_M2 0.018
r 50000_6000_M2 52000_6000_M2 0.018
r 52000_6000_M2 54000_6000_M2 0.018
r 54000_6000_M2 56000_6000_M2 0.018
r 56000_6000_M2 58000_6000_M2 0.018
r 58000_6000_M2 60000_6000_M2 0.018
r 60000_6000_M2 62000_6000_M2 0.018
r 62000_6000_M2 64000_6000_M2 0.018
r 64000_6000_M2 66000_6000_M2 0.018
r 66000_6000_M2 68000_6000_M2 0.018
r 68000_6000_M2 70000_6000_M2 0.018
r 70000_6000_M2 72000_6000_M2 0.018
r 72000_6000_M2 74000_6000_M2 0.018
r 74000_6000_M2 76000_6000_M2 0.018
r 76000_6000_M2 78000_6000_M2 0.018
r 78000_6000_M2 80000_6000_M2 0.018
r 80000_6000_M2 82000_6000_M2 0.018
r 82000_6000_M2 84000_6000_M2 0.018
r 84000_6000_M2 86000_6000_M2 0.018
r 86000_6000_M2 88000_6000_M2 0.018
r 88000_6000_M2 90000_6000_M2 0.018
r 90000_6000_M2 92000_6000_M2 0.018
r 92000_6000_M2 94000_6000_M2 0.018
r 94000_6000_M2 96000_6000_M2 0.018
r 96000_6000_M2 98000_6000_M2 0.018
r 98000_6000_M2 100000_6000_M2 0.018
r 2000_8000_M2 4000_8000_M2 0.018
r 4000_8000_M2 6000_8000_M2 0.018
r 6000_8000_M2 8000_8000_M2 0.018
r 8000_8000_M2 10000_8000_M2 0.018
r 10000_8000_M2 12000_8000_M2 0.018
r 12000_8000_M2 14000_8000_M2 0.018
r 14000_8000_M2 16000_8000_M2 0.018
r 16000_8000_M2 18000_8000_M2 0.018
r 18000_8000_M2 20000_8000_M2 0.018
r 20000_8000_M2 22000_8000_M2 0.018
r 22000_8000_M2 24000_8000_M2 0.018
r 24000_8000_M2 26000_8000_M2 0.018
r 26000_8000_M2 28000_8000_M2 0.018
r 28000_8000_M2 30000_8000_M2 0.018
r 30000_8000_M2 32000_8000_M2 0.018
r 32000_8000_M2 34000_8000_M2 0.018
r 34000_8000_M2 36000_8000_M2 0.018
r 36000_8000_M2 38000_8000_M2 0.018
r 38000_8000_M2 40000_8000_M2 0.018
r 40000_8000_M2 42000_8000_M2 0.018
r 42000_8000_M2 44000_8000_M2 0.018
r 44000_8000_M2 46000_8000_M2 0.018
r 46000_8000_M2 48000_8000_M2 0.018
r 48000_8000_M2 50000_8000_M2 0.018
r 50000_8000_M2 52000_8000_M2 0.018
r 52000_8000_M2 54000_8000_M2 0.018
r 54000_8000_M2 56000_8000_M2 0.018
r 56000_8000_M2 58000_8000_M2 0.018
r 58000_8000_M2 60000_8000_M2 0.018
r 60000_8000_M2 62000_8000_M2 0.018
r 62000_8000_M2 64000_8000_M2 0.018
r 64000_8000_M2 66000_8000_M2 0.018
r 66000_8000_M2 68000_8000_M2 0.018
r 68000_8000_M2 70000_8000_M2 0.018
r 70000_8000_M2 72000_8000_M2 0.018
r 72000_8000_M2 74000_8000_M2 0.018
r 74000_8000_M2 76000_8000_M2 0.018
r 76000_8000_M2 78000_8000_M2 0.018
r 78000_8000_M2 80000_8000_M2 0.018
r 80000_8000_M2 82000_8000_M2 0.018
r 82000_8000_M2 84000_8000_M2 0.018
r 84000_8000_M2 86000_8000_M2 0.018
r 86000_8000_M2 88000_8000_M2 0.018
r 88000_8000_M2 90000_8000_M2 0.018
r 90000_8000_M2 92000_8000_M2 0.018
r 92000_8000_M2 94000_8000_M2 0.018
r 94000_8000_M2 96000_8000_M2 0.018
r 96000_8000_M2 98000_8000_M2 0.018
r 98000_8000_M2 100000_8000_M2 0.018
r 2000_10000_M2 4000_10000_M2 0.018
r 4000_10000_M2 6000_10000_M2 0.018
r 6000_10000_M2 8000_10000_M2 0.018
r 8000_10000_M2 10000_10000_M2 0.018
r 10000_10000_M2 12000_10000_M2 0.018
r 12000_10000_M2 14000_10000_M2 0.018
r 14000_10000_M2 16000_10000_M2 0.018
r 16000_10000_M2 18000_10000_M2 0.018
r 18000_10000_M2 20000_10000_M2 0.018
r 20000_10000_M2 22000_10000_M2 0.018
r 22000_10000_M2 24000_10000_M2 0.018
r 24000_10000_M2 26000_10000_M2 0.018
r 26000_10000_M2 28000_10000_M2 0.018
r 28000_10000_M2 30000_10000_M2 0.018
r 30000_10000_M2 32000_10000_M2 0.018
r 32000_10000_M2 34000_10000_M2 0.018
r 34000_10000_M2 36000_10000_M2 0.018
r 36000_10000_M2 38000_10000_M2 0.018
r 38000_10000_M2 40000_10000_M2 0.018
r 40000_10000_M2 42000_10000_M2 0.018
r 42000_10000_M2 44000_10000_M2 0.018
r 44000_10000_M2 46000_10000_M2 0.018
r 46000_10000_M2 48000_10000_M2 0.018
r 48000_10000_M2 50000_10000_M2 0.018
r 50000_10000_M2 52000_10000_M2 0.018
r 52000_10000_M2 54000_10000_M2 0.018
r 54000_10000_M2 56000_10000_M2 0.018
r 56000_10000_M2 58000_10000_M2 0.018
r 58000_10000_M2 60000_10000_M2 0.018
r 60000_10000_M2 62000_10000_M2 0.018
r 62000_10000_M2 64000_10000_M2 0.018
r 64000_10000_M2 66000_10000_M2 0.018
r 66000_10000_M2 68000_10000_M2 0.018
r 68000_10000_M2 70000_10000_M2 0.018
r 70000_10000_M2 72000_10000_M2 0.018
r 72000_10000_M2 74000_10000_M2 0.018
r 74000_10000_M2 76000_10000_M2 0.018
r 76000_10000_M2 78000_10000_M2 0.018
r 78000_10000_M2 80000_10000_M2 0.018
r 80000_10000_M2 82000_10000_M2 0.018
r 82000_10000_M2 84000_10000_M2 0.018
r 84000_10000_M2 86000_10000_M2 0.018
r 86000_10000_M2 88000_10000_M2 0.018
r 88000_10000_M2 90000_10000_M2 0.018
r 90000_10000_M2 92000_10000_M2 0.018
r 92000_10000_M2 94000_10000_M2 0.018
r 94000_10000_M2 96000_10000_M2 0.018
r 96000_10000_M2 98000_10000_M2 0.018
r 98000_10000_M2 100000_10000_M2 0.018
r 2000_12000_M2 4000_12000_M2 0.018
r 4000_12000_M2 6000_12000_M2 0.018
r 6000_12000_M2 8000_12000_M2 0.018
r 8000_12000_M2 10000_12000_M2 0.018
r 10000_12000_M2 12000_12000_M2 0.018
r 12000_12000_M2 14000_12000_M2 0.018
r 14000_12000_M2 16000_12000_M2 0.018
r 16000_12000_M2 18000_12000_M2 0.018
r 18000_12000_M2 20000_12000_M2 0.018
r 20000_12000_M2 22000_12000_M2 0.018
r 22000_12000_M2 24000_12000_M2 0.018
r 24000_12000_M2 26000_12000_M2 0.018
r 26000_12000_M2 28000_12000_M2 0.018
r 28000_12000_M2 30000_12000_M2 0.018
r 30000_12000_M2 32000_12000_M2 0.018
r 32000_12000_M2 34000_12000_M2 0.018
r 34000_12000_M2 36000_12000_M2 0.018
r 36000_12000_M2 38000_12000_M2 0.018
r 38000_12000_M2 40000_12000_M2 0.018
r 40000_12000_M2 42000_12000_M2 0.018
r 42000_12000_M2 44000_12000_M2 0.018
r 44000_12000_M2 46000_12000_M2 0.018
r 46000_12000_M2 48000_12000_M2 0.018
r 48000_12000_M2 50000_12000_M2 0.018
r 50000_12000_M2 52000_12000_M2 0.018
r 52000_12000_M2 54000_12000_M2 0.018
r 54000_12000_M2 56000_12000_M2 0.018
r 56000_12000_M2 58000_12000_M2 0.018
r 58000_12000_M2 60000_12000_M2 0.018
r 60000_12000_M2 62000_12000_M2 0.018
r 62000_12000_M2 64000_12000_M2 0.018
r 64000_12000_M2 66000_12000_M2 0.018
r 66000_12000_M2 68000_12000_M2 0.018
r 68000_12000_M2 70000_12000_M2 0.018
r 70000_12000_M2 72000_12000_M2 0.018
r 72000_12000_M2 74000_12000_M2 0.018
r 74000_12000_M2 76000_12000_M2 0.018
r 76000_12000_M2 78000_12000_M2 0.018
r 78000_12000_M2 80000_12000_M2 0.018
r 80000_12000_M2 82000_12000_M2 0.018
r 82000_12000_M2 84000_12000_M2 0.018
r 84000_12000_M2 86000_12000_M2 0.018
r 86000_12000_M2 88000_12000_M2 0.018
r 88000_12000_M2 90000_12000_M2 0.018
r 90000_12000_M2 92000_12000_M2 0.018
r 92000_12000_M2 94000_12000_M2 0.018
r 94000_12000_M2 96000_12000_M2 0.018
r 96000_12000_M2 98000_12000_M2 0.018
r 98000_12000_M2 100000_12000_M2 0.018
r 2000_14000_M2 4000_14000_M2 0.018
r 4000_14000_M2 6000_14000_M2 0.018
r 6000_14000_M2 8000_14000_M2 0.018
r 8000_14000_M2 10000_14000_M2 0.018
r 10000_14000_M2 12000_14000_M2 0.018
r 12000_14000_M2 14000_14000_M2 0.018
r 14000_14000_M2 16000_14000_M2 0.018
r 16000_14000_M2 18000_14000_M2 0.018
r 18000_14000_M2 20000_14000_M2 0.018
r 20000_14000_M2 22000_14000_M2 0.018
r 22000_14000_M2 24000_14000_M2 0.018
r 24000_14000_M2 26000_14000_M2 0.018
r 26000_14000_M2 28000_14000_M2 0.018
r 28000_14000_M2 30000_14000_M2 0.018
r 30000_14000_M2 32000_14000_M2 0.018
r 32000_14000_M2 34000_14000_M2 0.018
r 34000_14000_M2 36000_14000_M2 0.018
r 36000_14000_M2 38000_14000_M2 0.018
r 38000_14000_M2 40000_14000_M2 0.018
r 40000_14000_M2 42000_14000_M2 0.018
r 42000_14000_M2 44000_14000_M2 0.018
r 44000_14000_M2 46000_14000_M2 0.018
r 46000_14000_M2 48000_14000_M2 0.018
r 48000_14000_M2 50000_14000_M2 0.018
r 50000_14000_M2 52000_14000_M2 0.018
r 52000_14000_M2 54000_14000_M2 0.018
r 54000_14000_M2 56000_14000_M2 0.018
r 56000_14000_M2 58000_14000_M2 0.018
r 58000_14000_M2 60000_14000_M2 0.018
r 60000_14000_M2 62000_14000_M2 0.018
r 62000_14000_M2 64000_14000_M2 0.018
r 64000_14000_M2 66000_14000_M2 0.018
r 66000_14000_M2 68000_14000_M2 0.018
r 68000_14000_M2 70000_14000_M2 0.018
r 70000_14000_M2 72000_14000_M2 0.018
r 72000_14000_M2 74000_14000_M2 0.018
r 74000_14000_M2 76000_14000_M2 0.018
r 76000_14000_M2 78000_14000_M2 0.018
r 78000_14000_M2 80000_14000_M2 0.018
r 80000_14000_M2 82000_14000_M2 0.018
r 82000_14000_M2 84000_14000_M2 0.018
r 84000_14000_M2 86000_14000_M2 0.018
r 86000_14000_M2 88000_14000_M2 0.018
r 88000_14000_M2 90000_14000_M2 0.018
r 90000_14000_M2 92000_14000_M2 0.018
r 92000_14000_M2 94000_14000_M2 0.018
r 94000_14000_M2 96000_14000_M2 0.018
r 96000_14000_M2 98000_14000_M2 0.018
r 98000_14000_M2 100000_14000_M2 0.018
r 2000_16000_M2 4000_16000_M2 0.018
r 4000_16000_M2 6000_16000_M2 0.018
r 6000_16000_M2 8000_16000_M2 0.018
r 8000_16000_M2 10000_16000_M2 0.018
r 10000_16000_M2 12000_16000_M2 0.018
r 12000_16000_M2 14000_16000_M2 0.018
r 14000_16000_M2 16000_16000_M2 0.018
r 16000_16000_M2 18000_16000_M2 0.018
r 18000_16000_M2 20000_16000_M2 0.018
r 20000_16000_M2 22000_16000_M2 0.018
r 22000_16000_M2 24000_16000_M2 0.018
r 24000_16000_M2 26000_16000_M2 0.018
r 26000_16000_M2 28000_16000_M2 0.018
r 28000_16000_M2 30000_16000_M2 0.018
r 30000_16000_M2 32000_16000_M2 0.018
r 32000_16000_M2 34000_16000_M2 0.018
r 34000_16000_M2 36000_16000_M2 0.018
r 36000_16000_M2 38000_16000_M2 0.018
r 38000_16000_M2 40000_16000_M2 0.018
r 40000_16000_M2 42000_16000_M2 0.018
r 42000_16000_M2 44000_16000_M2 0.018
r 44000_16000_M2 46000_16000_M2 0.018
r 46000_16000_M2 48000_16000_M2 0.018
r 48000_16000_M2 50000_16000_M2 0.018
r 50000_16000_M2 52000_16000_M2 0.018
r 52000_16000_M2 54000_16000_M2 0.018
r 54000_16000_M2 56000_16000_M2 0.018
r 56000_16000_M2 58000_16000_M2 0.018
r 58000_16000_M2 60000_16000_M2 0.018
r 60000_16000_M2 62000_16000_M2 0.018
r 62000_16000_M2 64000_16000_M2 0.018
r 64000_16000_M2 66000_16000_M2 0.018
r 66000_16000_M2 68000_16000_M2 0.018
r 68000_16000_M2 70000_16000_M2 0.018
r 70000_16000_M2 72000_16000_M2 0.018
r 72000_16000_M2 74000_16000_M2 0.018
r 74000_16000_M2 76000_16000_M2 0.018
r 76000_16000_M2 78000_16000_M2 0.018
r 78000_16000_M2 80000_16000_M2 0.018
r 80000_16000_M2 82000_16000_M2 0.018
r 82000_16000_M2 84000_16000_M2 0.018
r 84000_16000_M2 86000_16000_M2 0.018
r 86000_16000_M2 88000_16000_M2 0.018
r 88000_16000_M2 90000_16000_M2 0.018
r 90000_16000_M2 92000_16000_M2 0.018
r 92000_16000_M2 94000_16000_M2 0.018
r 94000_16000_M2 96000_16000_M2 0.018
r 96000_16000_M2 98000_16000_M2 0.018
r 98000_16000_M2 100000_16000_M2 0.018
r 2000_18000_M2 4000_18000_M2 0.018
r 4000_18000_M2 6000_18000_M2 0.018
r 6000_18000_M2 8000_18000_M2 0.018
r 8000_18000_M2 10000_18000_M2 0.018
r 10000_18000_M2 12000_18000_M2 0.018
r 12000_18000_M2 14000_18000_M2 0.018
r 14000_18000_M2 16000_18000_M2 0.018
r 16000_18000_M2 18000_18000_M2 0.018
r 18000_18000_M2 20000_18000_M2 0.018
r 20000_18000_M2 22000_18000_M2 0.018
r 22000_18000_M2 24000_18000_M2 0.018
r 24000_18000_M2 26000_18000_M2 0.018
r 26000_18000_M2 28000_18000_M2 0.018
r 28000_18000_M2 30000_18000_M2 0.018
r 30000_18000_M2 32000_18000_M2 0.018
r 32000_18000_M2 34000_18000_M2 0.018
r 34000_18000_M2 36000_18000_M2 0.018
r 36000_18000_M2 38000_18000_M2 0.018
r 38000_18000_M2 40000_18000_M2 0.018
r 40000_18000_M2 42000_18000_M2 0.018
r 42000_18000_M2 44000_18000_M2 0.018
r 44000_18000_M2 46000_18000_M2 0.018
r 46000_18000_M2 48000_18000_M2 0.018
r 48000_18000_M2 50000_18000_M2 0.018
r 50000_18000_M2 52000_18000_M2 0.018
r 52000_18000_M2 54000_18000_M2 0.018
r 54000_18000_M2 56000_18000_M2 0.018
r 56000_18000_M2 58000_18000_M2 0.018
r 58000_18000_M2 60000_18000_M2 0.018
r 60000_18000_M2 62000_18000_M2 0.018
r 62000_18000_M2 64000_18000_M2 0.018
r 64000_18000_M2 66000_18000_M2 0.018
r 66000_18000_M2 68000_18000_M2 0.018
r 68000_18000_M2 70000_18000_M2 0.018
r 70000_18000_M2 72000_18000_M2 0.018
r 72000_18000_M2 74000_18000_M2 0.018
r 74000_18000_M2 76000_18000_M2 0.018
r 76000_18000_M2 78000_18000_M2 0.018
r 78000_18000_M2 80000_18000_M2 0.018
r 80000_18000_M2 82000_18000_M2 0.018
r 82000_18000_M2 84000_18000_M2 0.018
r 84000_18000_M2 86000_18000_M2 0.018
r 86000_18000_M2 88000_18000_M2 0.018
r 88000_18000_M2 90000_18000_M2 0.018
r 90000_18000_M2 92000_18000_M2 0.018
r 92000_18000_M2 94000_18000_M2 0.018
r 94000_18000_M2 96000_18000_M2 0.018
r 96000_18000_M2 98000_18000_M2 0.018
r 98000_18000_M2 100000_18000_M2 0.018
r 2000_20000_M2 4000_20000_M2 0.018
r 4000_20000_M2 6000_20000_M2 0.018
r 6000_20000_M2 8000_20000_M2 0.018
r 8000_20000_M2 10000_20000_M2 0.018
r 10000_20000_M2 12000_20000_M2 0.018
r 12000_20000_M2 14000_20000_M2 0.018
r 14000_20000_M2 16000_20000_M2 0.018
r 16000_20000_M2 18000_20000_M2 0.018
r 18000_20000_M2 20000_20000_M2 0.018
r 20000_20000_M2 22000_20000_M2 0.018
r 22000_20000_M2 24000_20000_M2 0.018
r 24000_20000_M2 26000_20000_M2 0.018
r 26000_20000_M2 28000_20000_M2 0.018
r 28000_20000_M2 30000_20000_M2 0.018
r 30000_20000_M2 32000_20000_M2 0.018
r 32000_20000_M2 34000_20000_M2 0.018
r 34000_20000_M2 36000_20000_M2 0.018
r 36000_20000_M2 38000_20000_M2 0.018
r 38000_20000_M2 40000_20000_M2 0.018
r 40000_20000_M2 42000_20000_M2 0.018
r 42000_20000_M2 44000_20000_M2 0.018
r 44000_20000_M2 46000_20000_M2 0.018
r 46000_20000_M2 48000_20000_M2 0.018
r 48000_20000_M2 50000_20000_M2 0.018
r 50000_20000_M2 52000_20000_M2 0.018
r 52000_20000_M2 54000_20000_M2 0.018
r 54000_20000_M2 56000_20000_M2 0.018
r 56000_20000_M2 58000_20000_M2 0.018
r 58000_20000_M2 60000_20000_M2 0.018
r 60000_20000_M2 62000_20000_M2 0.018
r 62000_20000_M2 64000_20000_M2 0.018
r 64000_20000_M2 66000_20000_M2 0.018
r 66000_20000_M2 68000_20000_M2 0.018
r 68000_20000_M2 70000_20000_M2 0.018
r 70000_20000_M2 72000_20000_M2 0.018
r 72000_20000_M2 74000_20000_M2 0.018
r 74000_20000_M2 76000_20000_M2 0.018
r 76000_20000_M2 78000_20000_M2 0.018
r 78000_20000_M2 80000_20000_M2 0.018
r 80000_20000_M2 82000_20000_M2 0.018
r 82000_20000_M2 84000_20000_M2 0.018
r 84000_20000_M2 86000_20000_M2 0.018
r 86000_20000_M2 88000_20000_M2 0.018
r 88000_20000_M2 90000_20000_M2 0.018
r 90000_20000_M2 92000_20000_M2 0.018
r 92000_20000_M2 94000_20000_M2 0.018
r 94000_20000_M2 96000_20000_M2 0.018
r 96000_20000_M2 98000_20000_M2 0.018
r 98000_20000_M2 100000_20000_M2 0.018
r 2000_22000_M2 4000_22000_M2 0.018
r 4000_22000_M2 6000_22000_M2 0.018
r 6000_22000_M2 8000_22000_M2 0.018
r 8000_22000_M2 10000_22000_M2 0.018
r 10000_22000_M2 12000_22000_M2 0.018
r 12000_22000_M2 14000_22000_M2 0.018
r 14000_22000_M2 16000_22000_M2 0.018
r 16000_22000_M2 18000_22000_M2 0.018
r 18000_22000_M2 20000_22000_M2 0.018
r 20000_22000_M2 22000_22000_M2 0.018
r 22000_22000_M2 24000_22000_M2 0.018
r 24000_22000_M2 26000_22000_M2 0.018
r 26000_22000_M2 28000_22000_M2 0.018
r 28000_22000_M2 30000_22000_M2 0.018
r 30000_22000_M2 32000_22000_M2 0.018
r 32000_22000_M2 34000_22000_M2 0.018
r 34000_22000_M2 36000_22000_M2 0.018
r 36000_22000_M2 38000_22000_M2 0.018
r 38000_22000_M2 40000_22000_M2 0.018
r 40000_22000_M2 42000_22000_M2 0.018
r 42000_22000_M2 44000_22000_M2 0.018
r 44000_22000_M2 46000_22000_M2 0.018
r 46000_22000_M2 48000_22000_M2 0.018
r 48000_22000_M2 50000_22000_M2 0.018
r 50000_22000_M2 52000_22000_M2 0.018
r 52000_22000_M2 54000_22000_M2 0.018
r 54000_22000_M2 56000_22000_M2 0.018
r 56000_22000_M2 58000_22000_M2 0.018
r 58000_22000_M2 60000_22000_M2 0.018
r 60000_22000_M2 62000_22000_M2 0.018
r 62000_22000_M2 64000_22000_M2 0.018
r 64000_22000_M2 66000_22000_M2 0.018
r 66000_22000_M2 68000_22000_M2 0.018
r 68000_22000_M2 70000_22000_M2 0.018
r 70000_22000_M2 72000_22000_M2 0.018
r 72000_22000_M2 74000_22000_M2 0.018
r 74000_22000_M2 76000_22000_M2 0.018
r 76000_22000_M2 78000_22000_M2 0.018
r 78000_22000_M2 80000_22000_M2 0.018
r 80000_22000_M2 82000_22000_M2 0.018
r 82000_22000_M2 84000_22000_M2 0.018
r 84000_22000_M2 86000_22000_M2 0.018
r 86000_22000_M2 88000_22000_M2 0.018
r 88000_22000_M2 90000_22000_M2 0.018
r 90000_22000_M2 92000_22000_M2 0.018
r 92000_22000_M2 94000_22000_M2 0.018
r 94000_22000_M2 96000_22000_M2 0.018
r 96000_22000_M2 98000_22000_M2 0.018
r 98000_22000_M2 100000_22000_M2 0.018
r 2000_24000_M2 4000_24000_M2 0.018
r 4000_24000_M2 6000_24000_M2 0.018
r 6000_24000_M2 8000_24000_M2 0.018
r 8000_24000_M2 10000_24000_M2 0.018
r 10000_24000_M2 12000_24000_M2 0.018
r 12000_24000_M2 14000_24000_M2 0.018
r 14000_24000_M2 16000_24000_M2 0.018
r 16000_24000_M2 18000_24000_M2 0.018
r 18000_24000_M2 20000_24000_M2 0.018
r 20000_24000_M2 22000_24000_M2 0.018
r 22000_24000_M2 24000_24000_M2 0.018
r 24000_24000_M2 26000_24000_M2 0.018
r 26000_24000_M2 28000_24000_M2 0.018
r 28000_24000_M2 30000_24000_M2 0.018
r 30000_24000_M2 32000_24000_M2 0.018
r 32000_24000_M2 34000_24000_M2 0.018
r 34000_24000_M2 36000_24000_M2 0.018
r 36000_24000_M2 38000_24000_M2 0.018
r 38000_24000_M2 40000_24000_M2 0.018
r 40000_24000_M2 42000_24000_M2 0.018
r 42000_24000_M2 44000_24000_M2 0.018
r 44000_24000_M2 46000_24000_M2 0.018
r 46000_24000_M2 48000_24000_M2 0.018
r 48000_24000_M2 50000_24000_M2 0.018
r 50000_24000_M2 52000_24000_M2 0.018
r 52000_24000_M2 54000_24000_M2 0.018
r 54000_24000_M2 56000_24000_M2 0.018
r 56000_24000_M2 58000_24000_M2 0.018
r 58000_24000_M2 60000_24000_M2 0.018
r 60000_24000_M2 62000_24000_M2 0.018
r 62000_24000_M2 64000_24000_M2 0.018
r 64000_24000_M2 66000_24000_M2 0.018
r 66000_24000_M2 68000_24000_M2 0.018
r 68000_24000_M2 70000_24000_M2 0.018
r 70000_24000_M2 72000_24000_M2 0.018
r 72000_24000_M2 74000_24000_M2 0.018
r 74000_24000_M2 76000_24000_M2 0.018
r 76000_24000_M2 78000_24000_M2 0.018
r 78000_24000_M2 80000_24000_M2 0.018
r 80000_24000_M2 82000_24000_M2 0.018
r 82000_24000_M2 84000_24000_M2 0.018
r 84000_24000_M2 86000_24000_M2 0.018
r 86000_24000_M2 88000_24000_M2 0.018
r 88000_24000_M2 90000_24000_M2 0.018
r 90000_24000_M2 92000_24000_M2 0.018
r 92000_24000_M2 94000_24000_M2 0.018
r 94000_24000_M2 96000_24000_M2 0.018
r 96000_24000_M2 98000_24000_M2 0.018
r 98000_24000_M2 100000_24000_M2 0.018
r 2000_26000_M2 4000_26000_M2 0.018
r 4000_26000_M2 6000_26000_M2 0.018
r 6000_26000_M2 8000_26000_M2 0.018
r 8000_26000_M2 10000_26000_M2 0.018
r 10000_26000_M2 12000_26000_M2 0.018
r 12000_26000_M2 14000_26000_M2 0.018
r 14000_26000_M2 16000_26000_M2 0.018
r 16000_26000_M2 18000_26000_M2 0.018
r 18000_26000_M2 20000_26000_M2 0.018
r 20000_26000_M2 22000_26000_M2 0.018
r 22000_26000_M2 24000_26000_M2 0.018
r 24000_26000_M2 26000_26000_M2 0.018
r 26000_26000_M2 28000_26000_M2 0.018
r 28000_26000_M2 30000_26000_M2 0.018
r 30000_26000_M2 32000_26000_M2 0.018
r 32000_26000_M2 34000_26000_M2 0.018
r 34000_26000_M2 36000_26000_M2 0.018
r 36000_26000_M2 38000_26000_M2 0.018
r 38000_26000_M2 40000_26000_M2 0.018
r 40000_26000_M2 42000_26000_M2 0.018
r 42000_26000_M2 44000_26000_M2 0.018
r 44000_26000_M2 46000_26000_M2 0.018
r 46000_26000_M2 48000_26000_M2 0.018
r 48000_26000_M2 50000_26000_M2 0.018
r 50000_26000_M2 52000_26000_M2 0.018
r 52000_26000_M2 54000_26000_M2 0.018
r 54000_26000_M2 56000_26000_M2 0.018
r 56000_26000_M2 58000_26000_M2 0.018
r 58000_26000_M2 60000_26000_M2 0.018
r 60000_26000_M2 62000_26000_M2 0.018
r 62000_26000_M2 64000_26000_M2 0.018
r 64000_26000_M2 66000_26000_M2 0.018
r 66000_26000_M2 68000_26000_M2 0.018
r 68000_26000_M2 70000_26000_M2 0.018
r 70000_26000_M2 72000_26000_M2 0.018
r 72000_26000_M2 74000_26000_M2 0.018
r 74000_26000_M2 76000_26000_M2 0.018
r 76000_26000_M2 78000_26000_M2 0.018
r 78000_26000_M2 80000_26000_M2 0.018
r 80000_26000_M2 82000_26000_M2 0.018
r 82000_26000_M2 84000_26000_M2 0.018
r 84000_26000_M2 86000_26000_M2 0.018
r 86000_26000_M2 88000_26000_M2 0.018
r 88000_26000_M2 90000_26000_M2 0.018
r 90000_26000_M2 92000_26000_M2 0.018
r 92000_26000_M2 94000_26000_M2 0.018
r 94000_26000_M2 96000_26000_M2 0.018
r 96000_26000_M2 98000_26000_M2 0.018
r 98000_26000_M2 100000_26000_M2 0.018
r 2000_28000_M2 4000_28000_M2 0.018
r 4000_28000_M2 6000_28000_M2 0.018
r 6000_28000_M2 8000_28000_M2 0.018
r 8000_28000_M2 10000_28000_M2 0.018
r 10000_28000_M2 12000_28000_M2 0.018
r 12000_28000_M2 14000_28000_M2 0.018
r 14000_28000_M2 16000_28000_M2 0.018
r 16000_28000_M2 18000_28000_M2 0.018
r 18000_28000_M2 20000_28000_M2 0.018
r 20000_28000_M2 22000_28000_M2 0.018
r 22000_28000_M2 24000_28000_M2 0.018
r 24000_28000_M2 26000_28000_M2 0.018
r 26000_28000_M2 28000_28000_M2 0.018
r 28000_28000_M2 30000_28000_M2 0.018
r 30000_28000_M2 32000_28000_M2 0.018
r 32000_28000_M2 34000_28000_M2 0.018
r 34000_28000_M2 36000_28000_M2 0.018
r 36000_28000_M2 38000_28000_M2 0.018
r 38000_28000_M2 40000_28000_M2 0.018
r 40000_28000_M2 42000_28000_M2 0.018
r 42000_28000_M2 44000_28000_M2 0.018
r 44000_28000_M2 46000_28000_M2 0.018
r 46000_28000_M2 48000_28000_M2 0.018
r 48000_28000_M2 50000_28000_M2 0.018
r 50000_28000_M2 52000_28000_M2 0.018
r 52000_28000_M2 54000_28000_M2 0.018
r 54000_28000_M2 56000_28000_M2 0.018
r 56000_28000_M2 58000_28000_M2 0.018
r 58000_28000_M2 60000_28000_M2 0.018
r 60000_28000_M2 62000_28000_M2 0.018
r 62000_28000_M2 64000_28000_M2 0.018
r 64000_28000_M2 66000_28000_M2 0.018
r 66000_28000_M2 68000_28000_M2 0.018
r 68000_28000_M2 70000_28000_M2 0.018
r 70000_28000_M2 72000_28000_M2 0.018
r 72000_28000_M2 74000_28000_M2 0.018
r 74000_28000_M2 76000_28000_M2 0.018
r 76000_28000_M2 78000_28000_M2 0.018
r 78000_28000_M2 80000_28000_M2 0.018
r 80000_28000_M2 82000_28000_M2 0.018
r 82000_28000_M2 84000_28000_M2 0.018
r 84000_28000_M2 86000_28000_M2 0.018
r 86000_28000_M2 88000_28000_M2 0.018
r 88000_28000_M2 90000_28000_M2 0.018
r 90000_28000_M2 92000_28000_M2 0.018
r 92000_28000_M2 94000_28000_M2 0.018
r 94000_28000_M2 96000_28000_M2 0.018
r 96000_28000_M2 98000_28000_M2 0.018
r 98000_28000_M2 100000_28000_M2 0.018
r 2000_30000_M2 4000_30000_M2 0.018
r 4000_30000_M2 6000_30000_M2 0.018
r 6000_30000_M2 8000_30000_M2 0.018
r 8000_30000_M2 10000_30000_M2 0.018
r 10000_30000_M2 12000_30000_M2 0.018
r 12000_30000_M2 14000_30000_M2 0.018
r 14000_30000_M2 16000_30000_M2 0.018
r 16000_30000_M2 18000_30000_M2 0.018
r 18000_30000_M2 20000_30000_M2 0.018
r 20000_30000_M2 22000_30000_M2 0.018
r 22000_30000_M2 24000_30000_M2 0.018
r 24000_30000_M2 26000_30000_M2 0.018
r 26000_30000_M2 28000_30000_M2 0.018
r 28000_30000_M2 30000_30000_M2 0.018
r 30000_30000_M2 32000_30000_M2 0.018
r 32000_30000_M2 34000_30000_M2 0.018
r 34000_30000_M2 36000_30000_M2 0.018
r 36000_30000_M2 38000_30000_M2 0.018
r 38000_30000_M2 40000_30000_M2 0.018
r 40000_30000_M2 42000_30000_M2 0.018
r 42000_30000_M2 44000_30000_M2 0.018
r 44000_30000_M2 46000_30000_M2 0.018
r 46000_30000_M2 48000_30000_M2 0.018
r 48000_30000_M2 50000_30000_M2 0.018
r 50000_30000_M2 52000_30000_M2 0.018
r 52000_30000_M2 54000_30000_M2 0.018
r 54000_30000_M2 56000_30000_M2 0.018
r 56000_30000_M2 58000_30000_M2 0.018
r 58000_30000_M2 60000_30000_M2 0.018
r 60000_30000_M2 62000_30000_M2 0.018
r 62000_30000_M2 64000_30000_M2 0.018
r 64000_30000_M2 66000_30000_M2 0.018
r 66000_30000_M2 68000_30000_M2 0.018
r 68000_30000_M2 70000_30000_M2 0.018
r 70000_30000_M2 72000_30000_M2 0.018
r 72000_30000_M2 74000_30000_M2 0.018
r 74000_30000_M2 76000_30000_M2 0.018
r 76000_30000_M2 78000_30000_M2 0.018
r 78000_30000_M2 80000_30000_M2 0.018
r 80000_30000_M2 82000_30000_M2 0.018
r 82000_30000_M2 84000_30000_M2 0.018
r 84000_30000_M2 86000_30000_M2 0.018
r 86000_30000_M2 88000_30000_M2 0.018
r 88000_30000_M2 90000_30000_M2 0.018
r 90000_30000_M2 92000_30000_M2 0.018
r 92000_30000_M2 94000_30000_M2 0.018
r 94000_30000_M2 96000_30000_M2 0.018
r 96000_30000_M2 98000_30000_M2 0.018
r 98000_30000_M2 100000_30000_M2 0.018
r 2000_32000_M2 4000_32000_M2 0.018
r 4000_32000_M2 6000_32000_M2 0.018
r 6000_32000_M2 8000_32000_M2 0.018
r 8000_32000_M2 10000_32000_M2 0.018
r 10000_32000_M2 12000_32000_M2 0.018
r 12000_32000_M2 14000_32000_M2 0.018
r 14000_32000_M2 16000_32000_M2 0.018
r 16000_32000_M2 18000_32000_M2 0.018
r 18000_32000_M2 20000_32000_M2 0.018
r 20000_32000_M2 22000_32000_M2 0.018
r 22000_32000_M2 24000_32000_M2 0.018
r 24000_32000_M2 26000_32000_M2 0.018
r 26000_32000_M2 28000_32000_M2 0.018
r 28000_32000_M2 30000_32000_M2 0.018
r 30000_32000_M2 32000_32000_M2 0.018
r 32000_32000_M2 34000_32000_M2 0.018
r 34000_32000_M2 36000_32000_M2 0.018
r 36000_32000_M2 38000_32000_M2 0.018
r 38000_32000_M2 40000_32000_M2 0.018
r 40000_32000_M2 42000_32000_M2 0.018
r 42000_32000_M2 44000_32000_M2 0.018
r 44000_32000_M2 46000_32000_M2 0.018
r 46000_32000_M2 48000_32000_M2 0.018
r 48000_32000_M2 50000_32000_M2 0.018
r 50000_32000_M2 52000_32000_M2 0.018
r 52000_32000_M2 54000_32000_M2 0.018
r 54000_32000_M2 56000_32000_M2 0.018
r 56000_32000_M2 58000_32000_M2 0.018
r 58000_32000_M2 60000_32000_M2 0.018
r 60000_32000_M2 62000_32000_M2 0.018
r 62000_32000_M2 64000_32000_M2 0.018
r 64000_32000_M2 66000_32000_M2 0.018
r 66000_32000_M2 68000_32000_M2 0.018
r 68000_32000_M2 70000_32000_M2 0.018
r 70000_32000_M2 72000_32000_M2 0.018
r 72000_32000_M2 74000_32000_M2 0.018
r 74000_32000_M2 76000_32000_M2 0.018
r 76000_32000_M2 78000_32000_M2 0.018
r 78000_32000_M2 80000_32000_M2 0.018
r 80000_32000_M2 82000_32000_M2 0.018
r 82000_32000_M2 84000_32000_M2 0.018
r 84000_32000_M2 86000_32000_M2 0.018
r 86000_32000_M2 88000_32000_M2 0.018
r 88000_32000_M2 90000_32000_M2 0.018
r 90000_32000_M2 92000_32000_M2 0.018
r 92000_32000_M2 94000_32000_M2 0.018
r 94000_32000_M2 96000_32000_M2 0.018
r 96000_32000_M2 98000_32000_M2 0.018
r 98000_32000_M2 100000_32000_M2 0.018
r 2000_34000_M2 4000_34000_M2 0.018
r 4000_34000_M2 6000_34000_M2 0.018
r 6000_34000_M2 8000_34000_M2 0.018
r 8000_34000_M2 10000_34000_M2 0.018
r 10000_34000_M2 12000_34000_M2 0.018
r 12000_34000_M2 14000_34000_M2 0.018
r 14000_34000_M2 16000_34000_M2 0.018
r 16000_34000_M2 18000_34000_M2 0.018
r 18000_34000_M2 20000_34000_M2 0.018
r 20000_34000_M2 22000_34000_M2 0.018
r 22000_34000_M2 24000_34000_M2 0.018
r 24000_34000_M2 26000_34000_M2 0.018
r 26000_34000_M2 28000_34000_M2 0.018
r 28000_34000_M2 30000_34000_M2 0.018
r 30000_34000_M2 32000_34000_M2 0.018
r 32000_34000_M2 34000_34000_M2 0.018
r 34000_34000_M2 36000_34000_M2 0.018
r 36000_34000_M2 38000_34000_M2 0.018
r 38000_34000_M2 40000_34000_M2 0.018
r 40000_34000_M2 42000_34000_M2 0.018
r 42000_34000_M2 44000_34000_M2 0.018
r 44000_34000_M2 46000_34000_M2 0.018
r 46000_34000_M2 48000_34000_M2 0.018
r 48000_34000_M2 50000_34000_M2 0.018
r 50000_34000_M2 52000_34000_M2 0.018
r 52000_34000_M2 54000_34000_M2 0.018
r 54000_34000_M2 56000_34000_M2 0.018
r 56000_34000_M2 58000_34000_M2 0.018
r 58000_34000_M2 60000_34000_M2 0.018
r 60000_34000_M2 62000_34000_M2 0.018
r 62000_34000_M2 64000_34000_M2 0.018
r 64000_34000_M2 66000_34000_M2 0.018
r 66000_34000_M2 68000_34000_M2 0.018
r 68000_34000_M2 70000_34000_M2 0.018
r 70000_34000_M2 72000_34000_M2 0.018
r 72000_34000_M2 74000_34000_M2 0.018
r 74000_34000_M2 76000_34000_M2 0.018
r 76000_34000_M2 78000_34000_M2 0.018
r 78000_34000_M2 80000_34000_M2 0.018
r 80000_34000_M2 82000_34000_M2 0.018
r 82000_34000_M2 84000_34000_M2 0.018
r 84000_34000_M2 86000_34000_M2 0.018
r 86000_34000_M2 88000_34000_M2 0.018
r 88000_34000_M2 90000_34000_M2 0.018
r 90000_34000_M2 92000_34000_M2 0.018
r 92000_34000_M2 94000_34000_M2 0.018
r 94000_34000_M2 96000_34000_M2 0.018
r 96000_34000_M2 98000_34000_M2 0.018
r 98000_34000_M2 100000_34000_M2 0.018
r 2000_36000_M2 4000_36000_M2 0.018
r 4000_36000_M2 6000_36000_M2 0.018
r 6000_36000_M2 8000_36000_M2 0.018
r 8000_36000_M2 10000_36000_M2 0.018
r 10000_36000_M2 12000_36000_M2 0.018
r 12000_36000_M2 14000_36000_M2 0.018
r 14000_36000_M2 16000_36000_M2 0.018
r 16000_36000_M2 18000_36000_M2 0.018
r 18000_36000_M2 20000_36000_M2 0.018
r 20000_36000_M2 22000_36000_M2 0.018
r 22000_36000_M2 24000_36000_M2 0.018
r 24000_36000_M2 26000_36000_M2 0.018
r 26000_36000_M2 28000_36000_M2 0.018
r 28000_36000_M2 30000_36000_M2 0.018
r 30000_36000_M2 32000_36000_M2 0.018
r 32000_36000_M2 34000_36000_M2 0.018
r 34000_36000_M2 36000_36000_M2 0.018
r 36000_36000_M2 38000_36000_M2 0.018
r 38000_36000_M2 40000_36000_M2 0.018
r 40000_36000_M2 42000_36000_M2 0.018
r 42000_36000_M2 44000_36000_M2 0.018
r 44000_36000_M2 46000_36000_M2 0.018
r 46000_36000_M2 48000_36000_M2 0.018
r 48000_36000_M2 50000_36000_M2 0.018
r 50000_36000_M2 52000_36000_M2 0.018
r 52000_36000_M2 54000_36000_M2 0.018
r 54000_36000_M2 56000_36000_M2 0.018
r 56000_36000_M2 58000_36000_M2 0.018
r 58000_36000_M2 60000_36000_M2 0.018
r 60000_36000_M2 62000_36000_M2 0.018
r 62000_36000_M2 64000_36000_M2 0.018
r 64000_36000_M2 66000_36000_M2 0.018
r 66000_36000_M2 68000_36000_M2 0.018
r 68000_36000_M2 70000_36000_M2 0.018
r 70000_36000_M2 72000_36000_M2 0.018
r 72000_36000_M2 74000_36000_M2 0.018
r 74000_36000_M2 76000_36000_M2 0.018
r 76000_36000_M2 78000_36000_M2 0.018
r 78000_36000_M2 80000_36000_M2 0.018
r 80000_36000_M2 82000_36000_M2 0.018
r 82000_36000_M2 84000_36000_M2 0.018
r 84000_36000_M2 86000_36000_M2 0.018
r 86000_36000_M2 88000_36000_M2 0.018
r 88000_36000_M2 90000_36000_M2 0.018
r 90000_36000_M2 92000_36000_M2 0.018
r 92000_36000_M2 94000_36000_M2 0.018
r 94000_36000_M2 96000_36000_M2 0.018
r 96000_36000_M2 98000_36000_M2 0.018
r 98000_36000_M2 100000_36000_M2 0.018
r 2000_38000_M2 4000_38000_M2 0.018
r 4000_38000_M2 6000_38000_M2 0.018
r 6000_38000_M2 8000_38000_M2 0.018
r 8000_38000_M2 10000_38000_M2 0.018
r 10000_38000_M2 12000_38000_M2 0.018
r 12000_38000_M2 14000_38000_M2 0.018
r 14000_38000_M2 16000_38000_M2 0.018
r 16000_38000_M2 18000_38000_M2 0.018
r 18000_38000_M2 20000_38000_M2 0.018
r 20000_38000_M2 22000_38000_M2 0.018
r 22000_38000_M2 24000_38000_M2 0.018
r 24000_38000_M2 26000_38000_M2 0.018
r 26000_38000_M2 28000_38000_M2 0.018
r 28000_38000_M2 30000_38000_M2 0.018
r 30000_38000_M2 32000_38000_M2 0.018
r 32000_38000_M2 34000_38000_M2 0.018
r 34000_38000_M2 36000_38000_M2 0.018
r 36000_38000_M2 38000_38000_M2 0.018
r 38000_38000_M2 40000_38000_M2 0.018
r 40000_38000_M2 42000_38000_M2 0.018
r 42000_38000_M2 44000_38000_M2 0.018
r 44000_38000_M2 46000_38000_M2 0.018
r 46000_38000_M2 48000_38000_M2 0.018
r 48000_38000_M2 50000_38000_M2 0.018
r 50000_38000_M2 52000_38000_M2 0.018
r 52000_38000_M2 54000_38000_M2 0.018
r 54000_38000_M2 56000_38000_M2 0.018
r 56000_38000_M2 58000_38000_M2 0.018
r 58000_38000_M2 60000_38000_M2 0.018
r 60000_38000_M2 62000_38000_M2 0.018
r 62000_38000_M2 64000_38000_M2 0.018
r 64000_38000_M2 66000_38000_M2 0.018
r 66000_38000_M2 68000_38000_M2 0.018
r 68000_38000_M2 70000_38000_M2 0.018
r 70000_38000_M2 72000_38000_M2 0.018
r 72000_38000_M2 74000_38000_M2 0.018
r 74000_38000_M2 76000_38000_M2 0.018
r 76000_38000_M2 78000_38000_M2 0.018
r 78000_38000_M2 80000_38000_M2 0.018
r 80000_38000_M2 82000_38000_M2 0.018
r 82000_38000_M2 84000_38000_M2 0.018
r 84000_38000_M2 86000_38000_M2 0.018
r 86000_38000_M2 88000_38000_M2 0.018
r 88000_38000_M2 90000_38000_M2 0.018
r 90000_38000_M2 92000_38000_M2 0.018
r 92000_38000_M2 94000_38000_M2 0.018
r 94000_38000_M2 96000_38000_M2 0.018
r 96000_38000_M2 98000_38000_M2 0.018
r 98000_38000_M2 100000_38000_M2 0.018
r 2000_40000_M2 4000_40000_M2 0.018
r 4000_40000_M2 6000_40000_M2 0.018
r 6000_40000_M2 8000_40000_M2 0.018
r 8000_40000_M2 10000_40000_M2 0.018
r 10000_40000_M2 12000_40000_M2 0.018
r 12000_40000_M2 14000_40000_M2 0.018
r 14000_40000_M2 16000_40000_M2 0.018
r 16000_40000_M2 18000_40000_M2 0.018
r 18000_40000_M2 20000_40000_M2 0.018
r 20000_40000_M2 22000_40000_M2 0.018
r 22000_40000_M2 24000_40000_M2 0.018
r 24000_40000_M2 26000_40000_M2 0.018
r 26000_40000_M2 28000_40000_M2 0.018
r 28000_40000_M2 30000_40000_M2 0.018
r 30000_40000_M2 32000_40000_M2 0.018
r 32000_40000_M2 34000_40000_M2 0.018
r 34000_40000_M2 36000_40000_M2 0.018
r 36000_40000_M2 38000_40000_M2 0.018
r 38000_40000_M2 40000_40000_M2 0.018
r 40000_40000_M2 42000_40000_M2 0.018
r 42000_40000_M2 44000_40000_M2 0.018
r 44000_40000_M2 46000_40000_M2 0.018
r 46000_40000_M2 48000_40000_M2 0.018
r 48000_40000_M2 50000_40000_M2 0.018
r 50000_40000_M2 52000_40000_M2 0.018
r 52000_40000_M2 54000_40000_M2 0.018
r 54000_40000_M2 56000_40000_M2 0.018
r 56000_40000_M2 58000_40000_M2 0.018
r 58000_40000_M2 60000_40000_M2 0.018
r 60000_40000_M2 62000_40000_M2 0.018
r 62000_40000_M2 64000_40000_M2 0.018
r 64000_40000_M2 66000_40000_M2 0.018
r 66000_40000_M2 68000_40000_M2 0.018
r 68000_40000_M2 70000_40000_M2 0.018
r 70000_40000_M2 72000_40000_M2 0.018
r 72000_40000_M2 74000_40000_M2 0.018
r 74000_40000_M2 76000_40000_M2 0.018
r 76000_40000_M2 78000_40000_M2 0.018
r 78000_40000_M2 80000_40000_M2 0.018
r 80000_40000_M2 82000_40000_M2 0.018
r 82000_40000_M2 84000_40000_M2 0.018
r 84000_40000_M2 86000_40000_M2 0.018
r 86000_40000_M2 88000_40000_M2 0.018
r 88000_40000_M2 90000_40000_M2 0.018
r 90000_40000_M2 92000_40000_M2 0.018
r 92000_40000_M2 94000_40000_M2 0.018
r 94000_40000_M2 96000_40000_M2 0.018
r 96000_40000_M2 98000_40000_M2 0.018
r 98000_40000_M2 100000_40000_M2 0.018
r 2000_42000_M2 4000_42000_M2 0.018
r 4000_42000_M2 6000_42000_M2 0.018
r 6000_42000_M2 8000_42000_M2 0.018
r 8000_42000_M2 10000_42000_M2 0.018
r 10000_42000_M2 12000_42000_M2 0.018
r 12000_42000_M2 14000_42000_M2 0.018
r 14000_42000_M2 16000_42000_M2 0.018
r 16000_42000_M2 18000_42000_M2 0.018
r 18000_42000_M2 20000_42000_M2 0.018
r 20000_42000_M2 22000_42000_M2 0.018
r 22000_42000_M2 24000_42000_M2 0.018
r 24000_42000_M2 26000_42000_M2 0.018
r 26000_42000_M2 28000_42000_M2 0.018
r 28000_42000_M2 30000_42000_M2 0.018
r 30000_42000_M2 32000_42000_M2 0.018
r 32000_42000_M2 34000_42000_M2 0.018
r 34000_42000_M2 36000_42000_M2 0.018
r 36000_42000_M2 38000_42000_M2 0.018
r 38000_42000_M2 40000_42000_M2 0.018
r 40000_42000_M2 42000_42000_M2 0.018
r 42000_42000_M2 44000_42000_M2 0.018
r 44000_42000_M2 46000_42000_M2 0.018
r 46000_42000_M2 48000_42000_M2 0.018
r 48000_42000_M2 50000_42000_M2 0.018
r 50000_42000_M2 52000_42000_M2 0.018
r 52000_42000_M2 54000_42000_M2 0.018
r 54000_42000_M2 56000_42000_M2 0.018
r 56000_42000_M2 58000_42000_M2 0.018
r 58000_42000_M2 60000_42000_M2 0.018
r 60000_42000_M2 62000_42000_M2 0.018
r 62000_42000_M2 64000_42000_M2 0.018
r 64000_42000_M2 66000_42000_M2 0.018
r 66000_42000_M2 68000_42000_M2 0.018
r 68000_42000_M2 70000_42000_M2 0.018
r 70000_42000_M2 72000_42000_M2 0.018
r 72000_42000_M2 74000_42000_M2 0.018
r 74000_42000_M2 76000_42000_M2 0.018
r 76000_42000_M2 78000_42000_M2 0.018
r 78000_42000_M2 80000_42000_M2 0.018
r 80000_42000_M2 82000_42000_M2 0.018
r 82000_42000_M2 84000_42000_M2 0.018
r 84000_42000_M2 86000_42000_M2 0.018
r 86000_42000_M2 88000_42000_M2 0.018
r 88000_42000_M2 90000_42000_M2 0.018
r 90000_42000_M2 92000_42000_M2 0.018
r 92000_42000_M2 94000_42000_M2 0.018
r 94000_42000_M2 96000_42000_M2 0.018
r 96000_42000_M2 98000_42000_M2 0.018
r 98000_42000_M2 100000_42000_M2 0.018
r 2000_44000_M2 4000_44000_M2 0.018
r 4000_44000_M2 6000_44000_M2 0.018
r 6000_44000_M2 8000_44000_M2 0.018
r 8000_44000_M2 10000_44000_M2 0.018
r 10000_44000_M2 12000_44000_M2 0.018
r 12000_44000_M2 14000_44000_M2 0.018
r 14000_44000_M2 16000_44000_M2 0.018
r 16000_44000_M2 18000_44000_M2 0.018
r 18000_44000_M2 20000_44000_M2 0.018
r 20000_44000_M2 22000_44000_M2 0.018
r 22000_44000_M2 24000_44000_M2 0.018
r 24000_44000_M2 26000_44000_M2 0.018
r 26000_44000_M2 28000_44000_M2 0.018
r 28000_44000_M2 30000_44000_M2 0.018
r 30000_44000_M2 32000_44000_M2 0.018
r 32000_44000_M2 34000_44000_M2 0.018
r 34000_44000_M2 36000_44000_M2 0.018
r 36000_44000_M2 38000_44000_M2 0.018
r 38000_44000_M2 40000_44000_M2 0.018
r 40000_44000_M2 42000_44000_M2 0.018
r 42000_44000_M2 44000_44000_M2 0.018
r 44000_44000_M2 46000_44000_M2 0.018
r 46000_44000_M2 48000_44000_M2 0.018
r 48000_44000_M2 50000_44000_M2 0.018
r 50000_44000_M2 52000_44000_M2 0.018
r 52000_44000_M2 54000_44000_M2 0.018
r 54000_44000_M2 56000_44000_M2 0.018
r 56000_44000_M2 58000_44000_M2 0.018
r 58000_44000_M2 60000_44000_M2 0.018
r 60000_44000_M2 62000_44000_M2 0.018
r 62000_44000_M2 64000_44000_M2 0.018
r 64000_44000_M2 66000_44000_M2 0.018
r 66000_44000_M2 68000_44000_M2 0.018
r 68000_44000_M2 70000_44000_M2 0.018
r 70000_44000_M2 72000_44000_M2 0.018
r 72000_44000_M2 74000_44000_M2 0.018
r 74000_44000_M2 76000_44000_M2 0.018
r 76000_44000_M2 78000_44000_M2 0.018
r 78000_44000_M2 80000_44000_M2 0.018
r 80000_44000_M2 82000_44000_M2 0.018
r 82000_44000_M2 84000_44000_M2 0.018
r 84000_44000_M2 86000_44000_M2 0.018
r 86000_44000_M2 88000_44000_M2 0.018
r 88000_44000_M2 90000_44000_M2 0.018
r 90000_44000_M2 92000_44000_M2 0.018
r 92000_44000_M2 94000_44000_M2 0.018
r 94000_44000_M2 96000_44000_M2 0.018
r 96000_44000_M2 98000_44000_M2 0.018
r 98000_44000_M2 100000_44000_M2 0.018
r 2000_46000_M2 4000_46000_M2 0.018
r 4000_46000_M2 6000_46000_M2 0.018
r 6000_46000_M2 8000_46000_M2 0.018
r 8000_46000_M2 10000_46000_M2 0.018
r 10000_46000_M2 12000_46000_M2 0.018
r 12000_46000_M2 14000_46000_M2 0.018
r 14000_46000_M2 16000_46000_M2 0.018
r 16000_46000_M2 18000_46000_M2 0.018
r 18000_46000_M2 20000_46000_M2 0.018
r 20000_46000_M2 22000_46000_M2 0.018
r 22000_46000_M2 24000_46000_M2 0.018
r 24000_46000_M2 26000_46000_M2 0.018
r 26000_46000_M2 28000_46000_M2 0.018
r 28000_46000_M2 30000_46000_M2 0.018
r 30000_46000_M2 32000_46000_M2 0.018
r 32000_46000_M2 34000_46000_M2 0.018
r 34000_46000_M2 36000_46000_M2 0.018
r 36000_46000_M2 38000_46000_M2 0.018
r 38000_46000_M2 40000_46000_M2 0.018
r 40000_46000_M2 42000_46000_M2 0.018
r 42000_46000_M2 44000_46000_M2 0.018
r 44000_46000_M2 46000_46000_M2 0.018
r 46000_46000_M2 48000_46000_M2 0.018
r 48000_46000_M2 50000_46000_M2 0.018
r 50000_46000_M2 52000_46000_M2 0.018
r 52000_46000_M2 54000_46000_M2 0.018
r 54000_46000_M2 56000_46000_M2 0.018
r 56000_46000_M2 58000_46000_M2 0.018
r 58000_46000_M2 60000_46000_M2 0.018
r 60000_46000_M2 62000_46000_M2 0.018
r 62000_46000_M2 64000_46000_M2 0.018
r 64000_46000_M2 66000_46000_M2 0.018
r 66000_46000_M2 68000_46000_M2 0.018
r 68000_46000_M2 70000_46000_M2 0.018
r 70000_46000_M2 72000_46000_M2 0.018
r 72000_46000_M2 74000_46000_M2 0.018
r 74000_46000_M2 76000_46000_M2 0.018
r 76000_46000_M2 78000_46000_M2 0.018
r 78000_46000_M2 80000_46000_M2 0.018
r 80000_46000_M2 82000_46000_M2 0.018
r 82000_46000_M2 84000_46000_M2 0.018
r 84000_46000_M2 86000_46000_M2 0.018
r 86000_46000_M2 88000_46000_M2 0.018
r 88000_46000_M2 90000_46000_M2 0.018
r 90000_46000_M2 92000_46000_M2 0.018
r 92000_46000_M2 94000_46000_M2 0.018
r 94000_46000_M2 96000_46000_M2 0.018
r 96000_46000_M2 98000_46000_M2 0.018
r 98000_46000_M2 100000_46000_M2 0.018
r 2000_48000_M2 4000_48000_M2 0.018
r 4000_48000_M2 6000_48000_M2 0.018
r 6000_48000_M2 8000_48000_M2 0.018
r 8000_48000_M2 10000_48000_M2 0.018
r 10000_48000_M2 12000_48000_M2 0.018
r 12000_48000_M2 14000_48000_M2 0.018
r 14000_48000_M2 16000_48000_M2 0.018
r 16000_48000_M2 18000_48000_M2 0.018
r 18000_48000_M2 20000_48000_M2 0.018
r 20000_48000_M2 22000_48000_M2 0.018
r 22000_48000_M2 24000_48000_M2 0.018
r 24000_48000_M2 26000_48000_M2 0.018
r 26000_48000_M2 28000_48000_M2 0.018
r 28000_48000_M2 30000_48000_M2 0.018
r 30000_48000_M2 32000_48000_M2 0.018
r 32000_48000_M2 34000_48000_M2 0.018
r 34000_48000_M2 36000_48000_M2 0.018
r 36000_48000_M2 38000_48000_M2 0.018
r 38000_48000_M2 40000_48000_M2 0.018
r 40000_48000_M2 42000_48000_M2 0.018
r 42000_48000_M2 44000_48000_M2 0.018
r 44000_48000_M2 46000_48000_M2 0.018
r 46000_48000_M2 48000_48000_M2 0.018
r 48000_48000_M2 50000_48000_M2 0.018
r 50000_48000_M2 52000_48000_M2 0.018
r 52000_48000_M2 54000_48000_M2 0.018
r 54000_48000_M2 56000_48000_M2 0.018
r 56000_48000_M2 58000_48000_M2 0.018
r 58000_48000_M2 60000_48000_M2 0.018
r 60000_48000_M2 62000_48000_M2 0.018
r 62000_48000_M2 64000_48000_M2 0.018
r 64000_48000_M2 66000_48000_M2 0.018
r 66000_48000_M2 68000_48000_M2 0.018
r 68000_48000_M2 70000_48000_M2 0.018
r 70000_48000_M2 72000_48000_M2 0.018
r 72000_48000_M2 74000_48000_M2 0.018
r 74000_48000_M2 76000_48000_M2 0.018
r 76000_48000_M2 78000_48000_M2 0.018
r 78000_48000_M2 80000_48000_M2 0.018
r 80000_48000_M2 82000_48000_M2 0.018
r 82000_48000_M2 84000_48000_M2 0.018
r 84000_48000_M2 86000_48000_M2 0.018
r 86000_48000_M2 88000_48000_M2 0.018
r 88000_48000_M2 90000_48000_M2 0.018
r 90000_48000_M2 92000_48000_M2 0.018
r 92000_48000_M2 94000_48000_M2 0.018
r 94000_48000_M2 96000_48000_M2 0.018
r 96000_48000_M2 98000_48000_M2 0.018
r 98000_48000_M2 100000_48000_M2 0.018
r 2000_50000_M2 4000_50000_M2 0.018
r 4000_50000_M2 6000_50000_M2 0.018
r 6000_50000_M2 8000_50000_M2 0.018
r 8000_50000_M2 10000_50000_M2 0.018
r 10000_50000_M2 12000_50000_M2 0.018
r 12000_50000_M2 14000_50000_M2 0.018
r 14000_50000_M2 16000_50000_M2 0.018
r 16000_50000_M2 18000_50000_M2 0.018
r 18000_50000_M2 20000_50000_M2 0.018
r 20000_50000_M2 22000_50000_M2 0.018
r 22000_50000_M2 24000_50000_M2 0.018
r 24000_50000_M2 26000_50000_M2 0.018
r 26000_50000_M2 28000_50000_M2 0.018
r 28000_50000_M2 30000_50000_M2 0.018
r 30000_50000_M2 32000_50000_M2 0.018
r 32000_50000_M2 34000_50000_M2 0.018
r 34000_50000_M2 36000_50000_M2 0.018
r 36000_50000_M2 38000_50000_M2 0.018
r 38000_50000_M2 40000_50000_M2 0.018
r 40000_50000_M2 42000_50000_M2 0.018
r 42000_50000_M2 44000_50000_M2 0.018
r 44000_50000_M2 46000_50000_M2 0.018
r 46000_50000_M2 48000_50000_M2 0.018
r 48000_50000_M2 50000_50000_M2 0.018
r 50000_50000_M2 52000_50000_M2 0.018
r 52000_50000_M2 54000_50000_M2 0.018
r 54000_50000_M2 56000_50000_M2 0.018
r 56000_50000_M2 58000_50000_M2 0.018
r 58000_50000_M2 60000_50000_M2 0.018
r 60000_50000_M2 62000_50000_M2 0.018
r 62000_50000_M2 64000_50000_M2 0.018
r 64000_50000_M2 66000_50000_M2 0.018
r 66000_50000_M2 68000_50000_M2 0.018
r 68000_50000_M2 70000_50000_M2 0.018
r 70000_50000_M2 72000_50000_M2 0.018
r 72000_50000_M2 74000_50000_M2 0.018
r 74000_50000_M2 76000_50000_M2 0.018
r 76000_50000_M2 78000_50000_M2 0.018
r 78000_50000_M2 80000_50000_M2 0.018
r 80000_50000_M2 82000_50000_M2 0.018
r 82000_50000_M2 84000_50000_M2 0.018
r 84000_50000_M2 86000_50000_M2 0.018
r 86000_50000_M2 88000_50000_M2 0.018
r 88000_50000_M2 90000_50000_M2 0.018
r 90000_50000_M2 92000_50000_M2 0.018
r 92000_50000_M2 94000_50000_M2 0.018
r 94000_50000_M2 96000_50000_M2 0.018
r 96000_50000_M2 98000_50000_M2 0.018
r 98000_50000_M2 100000_50000_M2 0.018
r 2000_52000_M2 4000_52000_M2 0.018
r 4000_52000_M2 6000_52000_M2 0.018
r 6000_52000_M2 8000_52000_M2 0.018
r 8000_52000_M2 10000_52000_M2 0.018
r 10000_52000_M2 12000_52000_M2 0.018
r 12000_52000_M2 14000_52000_M2 0.018
r 14000_52000_M2 16000_52000_M2 0.018
r 16000_52000_M2 18000_52000_M2 0.018
r 18000_52000_M2 20000_52000_M2 0.018
r 20000_52000_M2 22000_52000_M2 0.018
r 22000_52000_M2 24000_52000_M2 0.018
r 24000_52000_M2 26000_52000_M2 0.018
r 26000_52000_M2 28000_52000_M2 0.018
r 28000_52000_M2 30000_52000_M2 0.018
r 30000_52000_M2 32000_52000_M2 0.018
r 32000_52000_M2 34000_52000_M2 0.018
r 34000_52000_M2 36000_52000_M2 0.018
r 36000_52000_M2 38000_52000_M2 0.018
r 38000_52000_M2 40000_52000_M2 0.018
r 40000_52000_M2 42000_52000_M2 0.018
r 42000_52000_M2 44000_52000_M2 0.018
r 44000_52000_M2 46000_52000_M2 0.018
r 46000_52000_M2 48000_52000_M2 0.018
r 48000_52000_M2 50000_52000_M2 0.018
r 50000_52000_M2 52000_52000_M2 0.018
r 52000_52000_M2 54000_52000_M2 0.018
r 54000_52000_M2 56000_52000_M2 0.018
r 56000_52000_M2 58000_52000_M2 0.018
r 58000_52000_M2 60000_52000_M2 0.018
r 60000_52000_M2 62000_52000_M2 0.018
r 62000_52000_M2 64000_52000_M2 0.018
r 64000_52000_M2 66000_52000_M2 0.018
r 66000_52000_M2 68000_52000_M2 0.018
r 68000_52000_M2 70000_52000_M2 0.018
r 70000_52000_M2 72000_52000_M2 0.018
r 72000_52000_M2 74000_52000_M2 0.018
r 74000_52000_M2 76000_52000_M2 0.018
r 76000_52000_M2 78000_52000_M2 0.018
r 78000_52000_M2 80000_52000_M2 0.018
r 80000_52000_M2 82000_52000_M2 0.018
r 82000_52000_M2 84000_52000_M2 0.018
r 84000_52000_M2 86000_52000_M2 0.018
r 86000_52000_M2 88000_52000_M2 0.018
r 88000_52000_M2 90000_52000_M2 0.018
r 90000_52000_M2 92000_52000_M2 0.018
r 92000_52000_M2 94000_52000_M2 0.018
r 94000_52000_M2 96000_52000_M2 0.018
r 96000_52000_M2 98000_52000_M2 0.018
r 98000_52000_M2 100000_52000_M2 0.018
r 2000_54000_M2 4000_54000_M2 0.018
r 4000_54000_M2 6000_54000_M2 0.018
r 6000_54000_M2 8000_54000_M2 0.018
r 8000_54000_M2 10000_54000_M2 0.018
r 10000_54000_M2 12000_54000_M2 0.018
r 12000_54000_M2 14000_54000_M2 0.018
r 14000_54000_M2 16000_54000_M2 0.018
r 16000_54000_M2 18000_54000_M2 0.018
r 18000_54000_M2 20000_54000_M2 0.018
r 20000_54000_M2 22000_54000_M2 0.018
r 22000_54000_M2 24000_54000_M2 0.018
r 24000_54000_M2 26000_54000_M2 0.018
r 26000_54000_M2 28000_54000_M2 0.018
r 28000_54000_M2 30000_54000_M2 0.018
r 30000_54000_M2 32000_54000_M2 0.018
r 32000_54000_M2 34000_54000_M2 0.018
r 34000_54000_M2 36000_54000_M2 0.018
r 36000_54000_M2 38000_54000_M2 0.018
r 38000_54000_M2 40000_54000_M2 0.018
r 40000_54000_M2 42000_54000_M2 0.018
r 42000_54000_M2 44000_54000_M2 0.018
r 44000_54000_M2 46000_54000_M2 0.018
r 46000_54000_M2 48000_54000_M2 0.018
r 48000_54000_M2 50000_54000_M2 0.018
r 50000_54000_M2 52000_54000_M2 0.018
r 52000_54000_M2 54000_54000_M2 0.018
r 54000_54000_M2 56000_54000_M2 0.018
r 56000_54000_M2 58000_54000_M2 0.018
r 58000_54000_M2 60000_54000_M2 0.018
r 60000_54000_M2 62000_54000_M2 0.018
r 62000_54000_M2 64000_54000_M2 0.018
r 64000_54000_M2 66000_54000_M2 0.018
r 66000_54000_M2 68000_54000_M2 0.018
r 68000_54000_M2 70000_54000_M2 0.018
r 70000_54000_M2 72000_54000_M2 0.018
r 72000_54000_M2 74000_54000_M2 0.018
r 74000_54000_M2 76000_54000_M2 0.018
r 76000_54000_M2 78000_54000_M2 0.018
r 78000_54000_M2 80000_54000_M2 0.018
r 80000_54000_M2 82000_54000_M2 0.018
r 82000_54000_M2 84000_54000_M2 0.018
r 84000_54000_M2 86000_54000_M2 0.018
r 86000_54000_M2 88000_54000_M2 0.018
r 88000_54000_M2 90000_54000_M2 0.018
r 90000_54000_M2 92000_54000_M2 0.018
r 92000_54000_M2 94000_54000_M2 0.018
r 94000_54000_M2 96000_54000_M2 0.018
r 96000_54000_M2 98000_54000_M2 0.018
r 98000_54000_M2 100000_54000_M2 0.018
r 2000_56000_M2 4000_56000_M2 0.018
r 4000_56000_M2 6000_56000_M2 0.018
r 6000_56000_M2 8000_56000_M2 0.018
r 8000_56000_M2 10000_56000_M2 0.018
r 10000_56000_M2 12000_56000_M2 0.018
r 12000_56000_M2 14000_56000_M2 0.018
r 14000_56000_M2 16000_56000_M2 0.018
r 16000_56000_M2 18000_56000_M2 0.018
r 18000_56000_M2 20000_56000_M2 0.018
r 20000_56000_M2 22000_56000_M2 0.018
r 22000_56000_M2 24000_56000_M2 0.018
r 24000_56000_M2 26000_56000_M2 0.018
r 26000_56000_M2 28000_56000_M2 0.018
r 28000_56000_M2 30000_56000_M2 0.018
r 30000_56000_M2 32000_56000_M2 0.018
r 32000_56000_M2 34000_56000_M2 0.018
r 34000_56000_M2 36000_56000_M2 0.018
r 36000_56000_M2 38000_56000_M2 0.018
r 38000_56000_M2 40000_56000_M2 0.018
r 40000_56000_M2 42000_56000_M2 0.018
r 42000_56000_M2 44000_56000_M2 0.018
r 44000_56000_M2 46000_56000_M2 0.018
r 46000_56000_M2 48000_56000_M2 0.018
r 48000_56000_M2 50000_56000_M2 0.018
r 50000_56000_M2 52000_56000_M2 0.018
r 52000_56000_M2 54000_56000_M2 0.018
r 54000_56000_M2 56000_56000_M2 0.018
r 56000_56000_M2 58000_56000_M2 0.018
r 58000_56000_M2 60000_56000_M2 0.018
r 60000_56000_M2 62000_56000_M2 0.018
r 62000_56000_M2 64000_56000_M2 0.018
r 64000_56000_M2 66000_56000_M2 0.018
r 66000_56000_M2 68000_56000_M2 0.018
r 68000_56000_M2 70000_56000_M2 0.018
r 70000_56000_M2 72000_56000_M2 0.018
r 72000_56000_M2 74000_56000_M2 0.018
r 74000_56000_M2 76000_56000_M2 0.018
r 76000_56000_M2 78000_56000_M2 0.018
r 78000_56000_M2 80000_56000_M2 0.018
r 80000_56000_M2 82000_56000_M2 0.018
r 82000_56000_M2 84000_56000_M2 0.018
r 84000_56000_M2 86000_56000_M2 0.018
r 86000_56000_M2 88000_56000_M2 0.018
r 88000_56000_M2 90000_56000_M2 0.018
r 90000_56000_M2 92000_56000_M2 0.018
r 92000_56000_M2 94000_56000_M2 0.018
r 94000_56000_M2 96000_56000_M2 0.018
r 96000_56000_M2 98000_56000_M2 0.018
r 98000_56000_M2 100000_56000_M2 0.018
r 2000_58000_M2 4000_58000_M2 0.018
r 4000_58000_M2 6000_58000_M2 0.018
r 6000_58000_M2 8000_58000_M2 0.018
r 8000_58000_M2 10000_58000_M2 0.018
r 10000_58000_M2 12000_58000_M2 0.018
r 12000_58000_M2 14000_58000_M2 0.018
r 14000_58000_M2 16000_58000_M2 0.018
r 16000_58000_M2 18000_58000_M2 0.018
r 18000_58000_M2 20000_58000_M2 0.018
r 20000_58000_M2 22000_58000_M2 0.018
r 22000_58000_M2 24000_58000_M2 0.018
r 24000_58000_M2 26000_58000_M2 0.018
r 26000_58000_M2 28000_58000_M2 0.018
r 28000_58000_M2 30000_58000_M2 0.018
r 30000_58000_M2 32000_58000_M2 0.018
r 32000_58000_M2 34000_58000_M2 0.018
r 34000_58000_M2 36000_58000_M2 0.018
r 36000_58000_M2 38000_58000_M2 0.018
r 38000_58000_M2 40000_58000_M2 0.018
r 40000_58000_M2 42000_58000_M2 0.018
r 42000_58000_M2 44000_58000_M2 0.018
r 44000_58000_M2 46000_58000_M2 0.018
r 46000_58000_M2 48000_58000_M2 0.018
r 48000_58000_M2 50000_58000_M2 0.018
r 50000_58000_M2 52000_58000_M2 0.018
r 52000_58000_M2 54000_58000_M2 0.018
r 54000_58000_M2 56000_58000_M2 0.018
r 56000_58000_M2 58000_58000_M2 0.018
r 58000_58000_M2 60000_58000_M2 0.018
r 60000_58000_M2 62000_58000_M2 0.018
r 62000_58000_M2 64000_58000_M2 0.018
r 64000_58000_M2 66000_58000_M2 0.018
r 66000_58000_M2 68000_58000_M2 0.018
r 68000_58000_M2 70000_58000_M2 0.018
r 70000_58000_M2 72000_58000_M2 0.018
r 72000_58000_M2 74000_58000_M2 0.018
r 74000_58000_M2 76000_58000_M2 0.018
r 76000_58000_M2 78000_58000_M2 0.018
r 78000_58000_M2 80000_58000_M2 0.018
r 80000_58000_M2 82000_58000_M2 0.018
r 82000_58000_M2 84000_58000_M2 0.018
r 84000_58000_M2 86000_58000_M2 0.018
r 86000_58000_M2 88000_58000_M2 0.018
r 88000_58000_M2 90000_58000_M2 0.018
r 90000_58000_M2 92000_58000_M2 0.018
r 92000_58000_M2 94000_58000_M2 0.018
r 94000_58000_M2 96000_58000_M2 0.018
r 96000_58000_M2 98000_58000_M2 0.018
r 98000_58000_M2 100000_58000_M2 0.018
r 2000_60000_M2 4000_60000_M2 0.018
r 4000_60000_M2 6000_60000_M2 0.018
r 6000_60000_M2 8000_60000_M2 0.018
r 8000_60000_M2 10000_60000_M2 0.018
r 10000_60000_M2 12000_60000_M2 0.018
r 12000_60000_M2 14000_60000_M2 0.018
r 14000_60000_M2 16000_60000_M2 0.018
r 16000_60000_M2 18000_60000_M2 0.018
r 18000_60000_M2 20000_60000_M2 0.018
r 20000_60000_M2 22000_60000_M2 0.018
r 22000_60000_M2 24000_60000_M2 0.018
r 24000_60000_M2 26000_60000_M2 0.018
r 26000_60000_M2 28000_60000_M2 0.018
r 28000_60000_M2 30000_60000_M2 0.018
r 30000_60000_M2 32000_60000_M2 0.018
r 32000_60000_M2 34000_60000_M2 0.018
r 34000_60000_M2 36000_60000_M2 0.018
r 36000_60000_M2 38000_60000_M2 0.018
r 38000_60000_M2 40000_60000_M2 0.018
r 40000_60000_M2 42000_60000_M2 0.018
r 42000_60000_M2 44000_60000_M2 0.018
r 44000_60000_M2 46000_60000_M2 0.018
r 46000_60000_M2 48000_60000_M2 0.018
r 48000_60000_M2 50000_60000_M2 0.018
r 50000_60000_M2 52000_60000_M2 0.018
r 52000_60000_M2 54000_60000_M2 0.018
r 54000_60000_M2 56000_60000_M2 0.018
r 56000_60000_M2 58000_60000_M2 0.018
r 58000_60000_M2 60000_60000_M2 0.018
r 60000_60000_M2 62000_60000_M2 0.018
r 62000_60000_M2 64000_60000_M2 0.018
r 64000_60000_M2 66000_60000_M2 0.018
r 66000_60000_M2 68000_60000_M2 0.018
r 68000_60000_M2 70000_60000_M2 0.018
r 70000_60000_M2 72000_60000_M2 0.018
r 72000_60000_M2 74000_60000_M2 0.018
r 74000_60000_M2 76000_60000_M2 0.018
r 76000_60000_M2 78000_60000_M2 0.018
r 78000_60000_M2 80000_60000_M2 0.018
r 80000_60000_M2 82000_60000_M2 0.018
r 82000_60000_M2 84000_60000_M2 0.018
r 84000_60000_M2 86000_60000_M2 0.018
r 86000_60000_M2 88000_60000_M2 0.018
r 88000_60000_M2 90000_60000_M2 0.018
r 90000_60000_M2 92000_60000_M2 0.018
r 92000_60000_M2 94000_60000_M2 0.018
r 94000_60000_M2 96000_60000_M2 0.018
r 96000_60000_M2 98000_60000_M2 0.018
r 98000_60000_M2 100000_60000_M2 0.018
r 2000_62000_M2 4000_62000_M2 0.018
r 4000_62000_M2 6000_62000_M2 0.018
r 6000_62000_M2 8000_62000_M2 0.018
r 8000_62000_M2 10000_62000_M2 0.018
r 10000_62000_M2 12000_62000_M2 0.018
r 12000_62000_M2 14000_62000_M2 0.018
r 14000_62000_M2 16000_62000_M2 0.018
r 16000_62000_M2 18000_62000_M2 0.018
r 18000_62000_M2 20000_62000_M2 0.018
r 20000_62000_M2 22000_62000_M2 0.018
r 22000_62000_M2 24000_62000_M2 0.018
r 24000_62000_M2 26000_62000_M2 0.018
r 26000_62000_M2 28000_62000_M2 0.018
r 28000_62000_M2 30000_62000_M2 0.018
r 30000_62000_M2 32000_62000_M2 0.018
r 32000_62000_M2 34000_62000_M2 0.018
r 34000_62000_M2 36000_62000_M2 0.018
r 36000_62000_M2 38000_62000_M2 0.018
r 38000_62000_M2 40000_62000_M2 0.018
r 40000_62000_M2 42000_62000_M2 0.018
r 42000_62000_M2 44000_62000_M2 0.018
r 44000_62000_M2 46000_62000_M2 0.018
r 46000_62000_M2 48000_62000_M2 0.018
r 48000_62000_M2 50000_62000_M2 0.018
r 50000_62000_M2 52000_62000_M2 0.018
r 52000_62000_M2 54000_62000_M2 0.018
r 54000_62000_M2 56000_62000_M2 0.018
r 56000_62000_M2 58000_62000_M2 0.018
r 58000_62000_M2 60000_62000_M2 0.018
r 60000_62000_M2 62000_62000_M2 0.018
r 62000_62000_M2 64000_62000_M2 0.018
r 64000_62000_M2 66000_62000_M2 0.018
r 66000_62000_M2 68000_62000_M2 0.018
r 68000_62000_M2 70000_62000_M2 0.018
r 70000_62000_M2 72000_62000_M2 0.018
r 72000_62000_M2 74000_62000_M2 0.018
r 74000_62000_M2 76000_62000_M2 0.018
r 76000_62000_M2 78000_62000_M2 0.018
r 78000_62000_M2 80000_62000_M2 0.018
r 80000_62000_M2 82000_62000_M2 0.018
r 82000_62000_M2 84000_62000_M2 0.018
r 84000_62000_M2 86000_62000_M2 0.018
r 86000_62000_M2 88000_62000_M2 0.018
r 88000_62000_M2 90000_62000_M2 0.018
r 90000_62000_M2 92000_62000_M2 0.018
r 92000_62000_M2 94000_62000_M2 0.018
r 94000_62000_M2 96000_62000_M2 0.018
r 96000_62000_M2 98000_62000_M2 0.018
r 98000_62000_M2 100000_62000_M2 0.018
r 2000_64000_M2 4000_64000_M2 0.018
r 4000_64000_M2 6000_64000_M2 0.018
r 6000_64000_M2 8000_64000_M2 0.018
r 8000_64000_M2 10000_64000_M2 0.018
r 10000_64000_M2 12000_64000_M2 0.018
r 12000_64000_M2 14000_64000_M2 0.018
r 14000_64000_M2 16000_64000_M2 0.018
r 16000_64000_M2 18000_64000_M2 0.018
r 18000_64000_M2 20000_64000_M2 0.018
r 20000_64000_M2 22000_64000_M2 0.018
r 22000_64000_M2 24000_64000_M2 0.018
r 24000_64000_M2 26000_64000_M2 0.018
r 26000_64000_M2 28000_64000_M2 0.018
r 28000_64000_M2 30000_64000_M2 0.018
r 30000_64000_M2 32000_64000_M2 0.018
r 32000_64000_M2 34000_64000_M2 0.018
r 34000_64000_M2 36000_64000_M2 0.018
r 36000_64000_M2 38000_64000_M2 0.018
r 38000_64000_M2 40000_64000_M2 0.018
r 40000_64000_M2 42000_64000_M2 0.018
r 42000_64000_M2 44000_64000_M2 0.018
r 44000_64000_M2 46000_64000_M2 0.018
r 46000_64000_M2 48000_64000_M2 0.018
r 48000_64000_M2 50000_64000_M2 0.018
r 50000_64000_M2 52000_64000_M2 0.018
r 52000_64000_M2 54000_64000_M2 0.018
r 54000_64000_M2 56000_64000_M2 0.018
r 56000_64000_M2 58000_64000_M2 0.018
r 58000_64000_M2 60000_64000_M2 0.018
r 60000_64000_M2 62000_64000_M2 0.018
r 62000_64000_M2 64000_64000_M2 0.018
r 64000_64000_M2 66000_64000_M2 0.018
r 66000_64000_M2 68000_64000_M2 0.018
r 68000_64000_M2 70000_64000_M2 0.018
r 70000_64000_M2 72000_64000_M2 0.018
r 72000_64000_M2 74000_64000_M2 0.018
r 74000_64000_M2 76000_64000_M2 0.018
r 76000_64000_M2 78000_64000_M2 0.018
r 78000_64000_M2 80000_64000_M2 0.018
r 80000_64000_M2 82000_64000_M2 0.018
r 82000_64000_M2 84000_64000_M2 0.018
r 84000_64000_M2 86000_64000_M2 0.018
r 86000_64000_M2 88000_64000_M2 0.018
r 88000_64000_M2 90000_64000_M2 0.018
r 90000_64000_M2 92000_64000_M2 0.018
r 92000_64000_M2 94000_64000_M2 0.018
r 94000_64000_M2 96000_64000_M2 0.018
r 96000_64000_M2 98000_64000_M2 0.018
r 98000_64000_M2 100000_64000_M2 0.018
r 2000_66000_M2 4000_66000_M2 0.018
r 4000_66000_M2 6000_66000_M2 0.018
r 6000_66000_M2 8000_66000_M2 0.018
r 8000_66000_M2 10000_66000_M2 0.018
r 10000_66000_M2 12000_66000_M2 0.018
r 12000_66000_M2 14000_66000_M2 0.018
r 14000_66000_M2 16000_66000_M2 0.018
r 16000_66000_M2 18000_66000_M2 0.018
r 18000_66000_M2 20000_66000_M2 0.018
r 20000_66000_M2 22000_66000_M2 0.018
r 22000_66000_M2 24000_66000_M2 0.018
r 24000_66000_M2 26000_66000_M2 0.018
r 26000_66000_M2 28000_66000_M2 0.018
r 28000_66000_M2 30000_66000_M2 0.018
r 30000_66000_M2 32000_66000_M2 0.018
r 32000_66000_M2 34000_66000_M2 0.018
r 34000_66000_M2 36000_66000_M2 0.018
r 36000_66000_M2 38000_66000_M2 0.018
r 38000_66000_M2 40000_66000_M2 0.018
r 40000_66000_M2 42000_66000_M2 0.018
r 42000_66000_M2 44000_66000_M2 0.018
r 44000_66000_M2 46000_66000_M2 0.018
r 46000_66000_M2 48000_66000_M2 0.018
r 48000_66000_M2 50000_66000_M2 0.018
r 50000_66000_M2 52000_66000_M2 0.018
r 52000_66000_M2 54000_66000_M2 0.018
r 54000_66000_M2 56000_66000_M2 0.018
r 56000_66000_M2 58000_66000_M2 0.018
r 58000_66000_M2 60000_66000_M2 0.018
r 60000_66000_M2 62000_66000_M2 0.018
r 62000_66000_M2 64000_66000_M2 0.018
r 64000_66000_M2 66000_66000_M2 0.018
r 66000_66000_M2 68000_66000_M2 0.018
r 68000_66000_M2 70000_66000_M2 0.018
r 70000_66000_M2 72000_66000_M2 0.018
r 72000_66000_M2 74000_66000_M2 0.018
r 74000_66000_M2 76000_66000_M2 0.018
r 76000_66000_M2 78000_66000_M2 0.018
r 78000_66000_M2 80000_66000_M2 0.018
r 80000_66000_M2 82000_66000_M2 0.018
r 82000_66000_M2 84000_66000_M2 0.018
r 84000_66000_M2 86000_66000_M2 0.018
r 86000_66000_M2 88000_66000_M2 0.018
r 88000_66000_M2 90000_66000_M2 0.018
r 90000_66000_M2 92000_66000_M2 0.018
r 92000_66000_M2 94000_66000_M2 0.018
r 94000_66000_M2 96000_66000_M2 0.018
r 96000_66000_M2 98000_66000_M2 0.018
r 98000_66000_M2 100000_66000_M2 0.018
r 2000_68000_M2 4000_68000_M2 0.018
r 4000_68000_M2 6000_68000_M2 0.018
r 6000_68000_M2 8000_68000_M2 0.018
r 8000_68000_M2 10000_68000_M2 0.018
r 10000_68000_M2 12000_68000_M2 0.018
r 12000_68000_M2 14000_68000_M2 0.018
r 14000_68000_M2 16000_68000_M2 0.018
r 16000_68000_M2 18000_68000_M2 0.018
r 18000_68000_M2 20000_68000_M2 0.018
r 20000_68000_M2 22000_68000_M2 0.018
r 22000_68000_M2 24000_68000_M2 0.018
r 24000_68000_M2 26000_68000_M2 0.018
r 26000_68000_M2 28000_68000_M2 0.018
r 28000_68000_M2 30000_68000_M2 0.018
r 30000_68000_M2 32000_68000_M2 0.018
r 32000_68000_M2 34000_68000_M2 0.018
r 34000_68000_M2 36000_68000_M2 0.018
r 36000_68000_M2 38000_68000_M2 0.018
r 38000_68000_M2 40000_68000_M2 0.018
r 40000_68000_M2 42000_68000_M2 0.018
r 42000_68000_M2 44000_68000_M2 0.018
r 44000_68000_M2 46000_68000_M2 0.018
r 46000_68000_M2 48000_68000_M2 0.018
r 48000_68000_M2 50000_68000_M2 0.018
r 50000_68000_M2 52000_68000_M2 0.018
r 52000_68000_M2 54000_68000_M2 0.018
r 54000_68000_M2 56000_68000_M2 0.018
r 56000_68000_M2 58000_68000_M2 0.018
r 58000_68000_M2 60000_68000_M2 0.018
r 60000_68000_M2 62000_68000_M2 0.018
r 62000_68000_M2 64000_68000_M2 0.018
r 64000_68000_M2 66000_68000_M2 0.018
r 66000_68000_M2 68000_68000_M2 0.018
r 68000_68000_M2 70000_68000_M2 0.018
r 70000_68000_M2 72000_68000_M2 0.018
r 72000_68000_M2 74000_68000_M2 0.018
r 74000_68000_M2 76000_68000_M2 0.018
r 76000_68000_M2 78000_68000_M2 0.018
r 78000_68000_M2 80000_68000_M2 0.018
r 80000_68000_M2 82000_68000_M2 0.018
r 82000_68000_M2 84000_68000_M2 0.018
r 84000_68000_M2 86000_68000_M2 0.018
r 86000_68000_M2 88000_68000_M2 0.018
r 88000_68000_M2 90000_68000_M2 0.018
r 90000_68000_M2 92000_68000_M2 0.018
r 92000_68000_M2 94000_68000_M2 0.018
r 94000_68000_M2 96000_68000_M2 0.018
r 96000_68000_M2 98000_68000_M2 0.018
r 98000_68000_M2 100000_68000_M2 0.018
r 2000_70000_M2 4000_70000_M2 0.018
r 4000_70000_M2 6000_70000_M2 0.018
r 6000_70000_M2 8000_70000_M2 0.018
r 8000_70000_M2 10000_70000_M2 0.018
r 10000_70000_M2 12000_70000_M2 0.018
r 12000_70000_M2 14000_70000_M2 0.018
r 14000_70000_M2 16000_70000_M2 0.018
r 16000_70000_M2 18000_70000_M2 0.018
r 18000_70000_M2 20000_70000_M2 0.018
r 20000_70000_M2 22000_70000_M2 0.018
r 22000_70000_M2 24000_70000_M2 0.018
r 24000_70000_M2 26000_70000_M2 0.018
r 26000_70000_M2 28000_70000_M2 0.018
r 28000_70000_M2 30000_70000_M2 0.018
r 30000_70000_M2 32000_70000_M2 0.018
r 32000_70000_M2 34000_70000_M2 0.018
r 34000_70000_M2 36000_70000_M2 0.018
r 36000_70000_M2 38000_70000_M2 0.018
r 38000_70000_M2 40000_70000_M2 0.018
r 40000_70000_M2 42000_70000_M2 0.018
r 42000_70000_M2 44000_70000_M2 0.018
r 44000_70000_M2 46000_70000_M2 0.018
r 46000_70000_M2 48000_70000_M2 0.018
r 48000_70000_M2 50000_70000_M2 0.018
r 50000_70000_M2 52000_70000_M2 0.018
r 52000_70000_M2 54000_70000_M2 0.018
r 54000_70000_M2 56000_70000_M2 0.018
r 56000_70000_M2 58000_70000_M2 0.018
r 58000_70000_M2 60000_70000_M2 0.018
r 60000_70000_M2 62000_70000_M2 0.018
r 62000_70000_M2 64000_70000_M2 0.018
r 64000_70000_M2 66000_70000_M2 0.018
r 66000_70000_M2 68000_70000_M2 0.018
r 68000_70000_M2 70000_70000_M2 0.018
r 70000_70000_M2 72000_70000_M2 0.018
r 72000_70000_M2 74000_70000_M2 0.018
r 74000_70000_M2 76000_70000_M2 0.018
r 76000_70000_M2 78000_70000_M2 0.018
r 78000_70000_M2 80000_70000_M2 0.018
r 80000_70000_M2 82000_70000_M2 0.018
r 82000_70000_M2 84000_70000_M2 0.018
r 84000_70000_M2 86000_70000_M2 0.018
r 86000_70000_M2 88000_70000_M2 0.018
r 88000_70000_M2 90000_70000_M2 0.018
r 90000_70000_M2 92000_70000_M2 0.018
r 92000_70000_M2 94000_70000_M2 0.018
r 94000_70000_M2 96000_70000_M2 0.018
r 96000_70000_M2 98000_70000_M2 0.018
r 98000_70000_M2 100000_70000_M2 0.018
r 2000_72000_M2 4000_72000_M2 0.018
r 4000_72000_M2 6000_72000_M2 0.018
r 6000_72000_M2 8000_72000_M2 0.018
r 8000_72000_M2 10000_72000_M2 0.018
r 10000_72000_M2 12000_72000_M2 0.018
r 12000_72000_M2 14000_72000_M2 0.018
r 14000_72000_M2 16000_72000_M2 0.018
r 16000_72000_M2 18000_72000_M2 0.018
r 18000_72000_M2 20000_72000_M2 0.018
r 20000_72000_M2 22000_72000_M2 0.018
r 22000_72000_M2 24000_72000_M2 0.018
r 24000_72000_M2 26000_72000_M2 0.018
r 26000_72000_M2 28000_72000_M2 0.018
r 28000_72000_M2 30000_72000_M2 0.018
r 30000_72000_M2 32000_72000_M2 0.018
r 32000_72000_M2 34000_72000_M2 0.018
r 34000_72000_M2 36000_72000_M2 0.018
r 36000_72000_M2 38000_72000_M2 0.018
r 38000_72000_M2 40000_72000_M2 0.018
r 40000_72000_M2 42000_72000_M2 0.018
r 42000_72000_M2 44000_72000_M2 0.018
r 44000_72000_M2 46000_72000_M2 0.018
r 46000_72000_M2 48000_72000_M2 0.018
r 48000_72000_M2 50000_72000_M2 0.018
r 50000_72000_M2 52000_72000_M2 0.018
r 52000_72000_M2 54000_72000_M2 0.018
r 54000_72000_M2 56000_72000_M2 0.018
r 56000_72000_M2 58000_72000_M2 0.018
r 58000_72000_M2 60000_72000_M2 0.018
r 60000_72000_M2 62000_72000_M2 0.018
r 62000_72000_M2 64000_72000_M2 0.018
r 64000_72000_M2 66000_72000_M2 0.018
r 66000_72000_M2 68000_72000_M2 0.018
r 68000_72000_M2 70000_72000_M2 0.018
r 70000_72000_M2 72000_72000_M2 0.018
r 72000_72000_M2 74000_72000_M2 0.018
r 74000_72000_M2 76000_72000_M2 0.018
r 76000_72000_M2 78000_72000_M2 0.018
r 78000_72000_M2 80000_72000_M2 0.018
r 80000_72000_M2 82000_72000_M2 0.018
r 82000_72000_M2 84000_72000_M2 0.018
r 84000_72000_M2 86000_72000_M2 0.018
r 86000_72000_M2 88000_72000_M2 0.018
r 88000_72000_M2 90000_72000_M2 0.018
r 90000_72000_M2 92000_72000_M2 0.018
r 92000_72000_M2 94000_72000_M2 0.018
r 94000_72000_M2 96000_72000_M2 0.018
r 96000_72000_M2 98000_72000_M2 0.018
r 98000_72000_M2 100000_72000_M2 0.018
r 2000_74000_M2 4000_74000_M2 0.018
r 4000_74000_M2 6000_74000_M2 0.018
r 6000_74000_M2 8000_74000_M2 0.018
r 8000_74000_M2 10000_74000_M2 0.018
r 10000_74000_M2 12000_74000_M2 0.018
r 12000_74000_M2 14000_74000_M2 0.018
r 14000_74000_M2 16000_74000_M2 0.018
r 16000_74000_M2 18000_74000_M2 0.018
r 18000_74000_M2 20000_74000_M2 0.018
r 20000_74000_M2 22000_74000_M2 0.018
r 22000_74000_M2 24000_74000_M2 0.018
r 24000_74000_M2 26000_74000_M2 0.018
r 26000_74000_M2 28000_74000_M2 0.018
r 28000_74000_M2 30000_74000_M2 0.018
r 30000_74000_M2 32000_74000_M2 0.018
r 32000_74000_M2 34000_74000_M2 0.018
r 34000_74000_M2 36000_74000_M2 0.018
r 36000_74000_M2 38000_74000_M2 0.018
r 38000_74000_M2 40000_74000_M2 0.018
r 40000_74000_M2 42000_74000_M2 0.018
r 42000_74000_M2 44000_74000_M2 0.018
r 44000_74000_M2 46000_74000_M2 0.018
r 46000_74000_M2 48000_74000_M2 0.018
r 48000_74000_M2 50000_74000_M2 0.018
r 50000_74000_M2 52000_74000_M2 0.018
r 52000_74000_M2 54000_74000_M2 0.018
r 54000_74000_M2 56000_74000_M2 0.018
r 56000_74000_M2 58000_74000_M2 0.018
r 58000_74000_M2 60000_74000_M2 0.018
r 60000_74000_M2 62000_74000_M2 0.018
r 62000_74000_M2 64000_74000_M2 0.018
r 64000_74000_M2 66000_74000_M2 0.018
r 66000_74000_M2 68000_74000_M2 0.018
r 68000_74000_M2 70000_74000_M2 0.018
r 70000_74000_M2 72000_74000_M2 0.018
r 72000_74000_M2 74000_74000_M2 0.018
r 74000_74000_M2 76000_74000_M2 0.018
r 76000_74000_M2 78000_74000_M2 0.018
r 78000_74000_M2 80000_74000_M2 0.018
r 80000_74000_M2 82000_74000_M2 0.018
r 82000_74000_M2 84000_74000_M2 0.018
r 84000_74000_M2 86000_74000_M2 0.018
r 86000_74000_M2 88000_74000_M2 0.018
r 88000_74000_M2 90000_74000_M2 0.018
r 90000_74000_M2 92000_74000_M2 0.018
r 92000_74000_M2 94000_74000_M2 0.018
r 94000_74000_M2 96000_74000_M2 0.018
r 96000_74000_M2 98000_74000_M2 0.018
r 98000_74000_M2 100000_74000_M2 0.018
r 2000_76000_M2 4000_76000_M2 0.018
r 4000_76000_M2 6000_76000_M2 0.018
r 6000_76000_M2 8000_76000_M2 0.018
r 8000_76000_M2 10000_76000_M2 0.018
r 10000_76000_M2 12000_76000_M2 0.018
r 12000_76000_M2 14000_76000_M2 0.018
r 14000_76000_M2 16000_76000_M2 0.018
r 16000_76000_M2 18000_76000_M2 0.018
r 18000_76000_M2 20000_76000_M2 0.018
r 20000_76000_M2 22000_76000_M2 0.018
r 22000_76000_M2 24000_76000_M2 0.018
r 24000_76000_M2 26000_76000_M2 0.018
r 26000_76000_M2 28000_76000_M2 0.018
r 28000_76000_M2 30000_76000_M2 0.018
r 30000_76000_M2 32000_76000_M2 0.018
r 32000_76000_M2 34000_76000_M2 0.018
r 34000_76000_M2 36000_76000_M2 0.018
r 36000_76000_M2 38000_76000_M2 0.018
r 38000_76000_M2 40000_76000_M2 0.018
r 40000_76000_M2 42000_76000_M2 0.018
r 42000_76000_M2 44000_76000_M2 0.018
r 44000_76000_M2 46000_76000_M2 0.018
r 46000_76000_M2 48000_76000_M2 0.018
r 48000_76000_M2 50000_76000_M2 0.018
r 50000_76000_M2 52000_76000_M2 0.018
r 52000_76000_M2 54000_76000_M2 0.018
r 54000_76000_M2 56000_76000_M2 0.018
r 56000_76000_M2 58000_76000_M2 0.018
r 58000_76000_M2 60000_76000_M2 0.018
r 60000_76000_M2 62000_76000_M2 0.018
r 62000_76000_M2 64000_76000_M2 0.018
r 64000_76000_M2 66000_76000_M2 0.018
r 66000_76000_M2 68000_76000_M2 0.018
r 68000_76000_M2 70000_76000_M2 0.018
r 70000_76000_M2 72000_76000_M2 0.018
r 72000_76000_M2 74000_76000_M2 0.018
r 74000_76000_M2 76000_76000_M2 0.018
r 76000_76000_M2 78000_76000_M2 0.018
r 78000_76000_M2 80000_76000_M2 0.018
r 80000_76000_M2 82000_76000_M2 0.018
r 82000_76000_M2 84000_76000_M2 0.018
r 84000_76000_M2 86000_76000_M2 0.018
r 86000_76000_M2 88000_76000_M2 0.018
r 88000_76000_M2 90000_76000_M2 0.018
r 90000_76000_M2 92000_76000_M2 0.018
r 92000_76000_M2 94000_76000_M2 0.018
r 94000_76000_M2 96000_76000_M2 0.018
r 96000_76000_M2 98000_76000_M2 0.018
r 98000_76000_M2 100000_76000_M2 0.018
r 2000_78000_M2 4000_78000_M2 0.018
r 4000_78000_M2 6000_78000_M2 0.018
r 6000_78000_M2 8000_78000_M2 0.018
r 8000_78000_M2 10000_78000_M2 0.018
r 10000_78000_M2 12000_78000_M2 0.018
r 12000_78000_M2 14000_78000_M2 0.018
r 14000_78000_M2 16000_78000_M2 0.018
r 16000_78000_M2 18000_78000_M2 0.018
r 18000_78000_M2 20000_78000_M2 0.018
r 20000_78000_M2 22000_78000_M2 0.018
r 22000_78000_M2 24000_78000_M2 0.018
r 24000_78000_M2 26000_78000_M2 0.018
r 26000_78000_M2 28000_78000_M2 0.018
r 28000_78000_M2 30000_78000_M2 0.018
r 30000_78000_M2 32000_78000_M2 0.018
r 32000_78000_M2 34000_78000_M2 0.018
r 34000_78000_M2 36000_78000_M2 0.018
r 36000_78000_M2 38000_78000_M2 0.018
r 38000_78000_M2 40000_78000_M2 0.018
r 40000_78000_M2 42000_78000_M2 0.018
r 42000_78000_M2 44000_78000_M2 0.018
r 44000_78000_M2 46000_78000_M2 0.018
r 46000_78000_M2 48000_78000_M2 0.018
r 48000_78000_M2 50000_78000_M2 0.018
r 50000_78000_M2 52000_78000_M2 0.018
r 52000_78000_M2 54000_78000_M2 0.018
r 54000_78000_M2 56000_78000_M2 0.018
r 56000_78000_M2 58000_78000_M2 0.018
r 58000_78000_M2 60000_78000_M2 0.018
r 60000_78000_M2 62000_78000_M2 0.018
r 62000_78000_M2 64000_78000_M2 0.018
r 64000_78000_M2 66000_78000_M2 0.018
r 66000_78000_M2 68000_78000_M2 0.018
r 68000_78000_M2 70000_78000_M2 0.018
r 70000_78000_M2 72000_78000_M2 0.018
r 72000_78000_M2 74000_78000_M2 0.018
r 74000_78000_M2 76000_78000_M2 0.018
r 76000_78000_M2 78000_78000_M2 0.018
r 78000_78000_M2 80000_78000_M2 0.018
r 80000_78000_M2 82000_78000_M2 0.018
r 82000_78000_M2 84000_78000_M2 0.018
r 84000_78000_M2 86000_78000_M2 0.018
r 86000_78000_M2 88000_78000_M2 0.018
r 88000_78000_M2 90000_78000_M2 0.018
r 90000_78000_M2 92000_78000_M2 0.018
r 92000_78000_M2 94000_78000_M2 0.018
r 94000_78000_M2 96000_78000_M2 0.018
r 96000_78000_M2 98000_78000_M2 0.018
r 98000_78000_M2 100000_78000_M2 0.018
r 2000_80000_M2 4000_80000_M2 0.018
r 4000_80000_M2 6000_80000_M2 0.018
r 6000_80000_M2 8000_80000_M2 0.018
r 8000_80000_M2 10000_80000_M2 0.018
r 10000_80000_M2 12000_80000_M2 0.018
r 12000_80000_M2 14000_80000_M2 0.018
r 14000_80000_M2 16000_80000_M2 0.018
r 16000_80000_M2 18000_80000_M2 0.018
r 18000_80000_M2 20000_80000_M2 0.018
r 20000_80000_M2 22000_80000_M2 0.018
r 22000_80000_M2 24000_80000_M2 0.018
r 24000_80000_M2 26000_80000_M2 0.018
r 26000_80000_M2 28000_80000_M2 0.018
r 28000_80000_M2 30000_80000_M2 0.018
r 30000_80000_M2 32000_80000_M2 0.018
r 32000_80000_M2 34000_80000_M2 0.018
r 34000_80000_M2 36000_80000_M2 0.018
r 36000_80000_M2 38000_80000_M2 0.018
r 38000_80000_M2 40000_80000_M2 0.018
r 40000_80000_M2 42000_80000_M2 0.018
r 42000_80000_M2 44000_80000_M2 0.018
r 44000_80000_M2 46000_80000_M2 0.018
r 46000_80000_M2 48000_80000_M2 0.018
r 48000_80000_M2 50000_80000_M2 0.018
r 50000_80000_M2 52000_80000_M2 0.018
r 52000_80000_M2 54000_80000_M2 0.018
r 54000_80000_M2 56000_80000_M2 0.018
r 56000_80000_M2 58000_80000_M2 0.018
r 58000_80000_M2 60000_80000_M2 0.018
r 60000_80000_M2 62000_80000_M2 0.018
r 62000_80000_M2 64000_80000_M2 0.018
r 64000_80000_M2 66000_80000_M2 0.018
r 66000_80000_M2 68000_80000_M2 0.018
r 68000_80000_M2 70000_80000_M2 0.018
r 70000_80000_M2 72000_80000_M2 0.018
r 72000_80000_M2 74000_80000_M2 0.018
r 74000_80000_M2 76000_80000_M2 0.018
r 76000_80000_M2 78000_80000_M2 0.018
r 78000_80000_M2 80000_80000_M2 0.018
r 80000_80000_M2 82000_80000_M2 0.018
r 82000_80000_M2 84000_80000_M2 0.018
r 84000_80000_M2 86000_80000_M2 0.018
r 86000_80000_M2 88000_80000_M2 0.018
r 88000_80000_M2 90000_80000_M2 0.018
r 90000_80000_M2 92000_80000_M2 0.018
r 92000_80000_M2 94000_80000_M2 0.018
r 94000_80000_M2 96000_80000_M2 0.018
r 96000_80000_M2 98000_80000_M2 0.018
r 98000_80000_M2 100000_80000_M2 0.018
r 2000_82000_M2 4000_82000_M2 0.018
r 4000_82000_M2 6000_82000_M2 0.018
r 6000_82000_M2 8000_82000_M2 0.018
r 8000_82000_M2 10000_82000_M2 0.018
r 10000_82000_M2 12000_82000_M2 0.018
r 12000_82000_M2 14000_82000_M2 0.018
r 14000_82000_M2 16000_82000_M2 0.018
r 16000_82000_M2 18000_82000_M2 0.018
r 18000_82000_M2 20000_82000_M2 0.018
r 20000_82000_M2 22000_82000_M2 0.018
r 22000_82000_M2 24000_82000_M2 0.018
r 24000_82000_M2 26000_82000_M2 0.018
r 26000_82000_M2 28000_82000_M2 0.018
r 28000_82000_M2 30000_82000_M2 0.018
r 30000_82000_M2 32000_82000_M2 0.018
r 32000_82000_M2 34000_82000_M2 0.018
r 34000_82000_M2 36000_82000_M2 0.018
r 36000_82000_M2 38000_82000_M2 0.018
r 38000_82000_M2 40000_82000_M2 0.018
r 40000_82000_M2 42000_82000_M2 0.018
r 42000_82000_M2 44000_82000_M2 0.018
r 44000_82000_M2 46000_82000_M2 0.018
r 46000_82000_M2 48000_82000_M2 0.018
r 48000_82000_M2 50000_82000_M2 0.018
r 50000_82000_M2 52000_82000_M2 0.018
r 52000_82000_M2 54000_82000_M2 0.018
r 54000_82000_M2 56000_82000_M2 0.018
r 56000_82000_M2 58000_82000_M2 0.018
r 58000_82000_M2 60000_82000_M2 0.018
r 60000_82000_M2 62000_82000_M2 0.018
r 62000_82000_M2 64000_82000_M2 0.018
r 64000_82000_M2 66000_82000_M2 0.018
r 66000_82000_M2 68000_82000_M2 0.018
r 68000_82000_M2 70000_82000_M2 0.018
r 70000_82000_M2 72000_82000_M2 0.018
r 72000_82000_M2 74000_82000_M2 0.018
r 74000_82000_M2 76000_82000_M2 0.018
r 76000_82000_M2 78000_82000_M2 0.018
r 78000_82000_M2 80000_82000_M2 0.018
r 80000_82000_M2 82000_82000_M2 0.018
r 82000_82000_M2 84000_82000_M2 0.018
r 84000_82000_M2 86000_82000_M2 0.018
r 86000_82000_M2 88000_82000_M2 0.018
r 88000_82000_M2 90000_82000_M2 0.018
r 90000_82000_M2 92000_82000_M2 0.018
r 92000_82000_M2 94000_82000_M2 0.018
r 94000_82000_M2 96000_82000_M2 0.018
r 96000_82000_M2 98000_82000_M2 0.018
r 98000_82000_M2 100000_82000_M2 0.018
r 2000_84000_M2 4000_84000_M2 0.018
r 4000_84000_M2 6000_84000_M2 0.018
r 6000_84000_M2 8000_84000_M2 0.018
r 8000_84000_M2 10000_84000_M2 0.018
r 10000_84000_M2 12000_84000_M2 0.018
r 12000_84000_M2 14000_84000_M2 0.018
r 14000_84000_M2 16000_84000_M2 0.018
r 16000_84000_M2 18000_84000_M2 0.018
r 18000_84000_M2 20000_84000_M2 0.018
r 20000_84000_M2 22000_84000_M2 0.018
r 22000_84000_M2 24000_84000_M2 0.018
r 24000_84000_M2 26000_84000_M2 0.018
r 26000_84000_M2 28000_84000_M2 0.018
r 28000_84000_M2 30000_84000_M2 0.018
r 30000_84000_M2 32000_84000_M2 0.018
r 32000_84000_M2 34000_84000_M2 0.018
r 34000_84000_M2 36000_84000_M2 0.018
r 36000_84000_M2 38000_84000_M2 0.018
r 38000_84000_M2 40000_84000_M2 0.018
r 40000_84000_M2 42000_84000_M2 0.018
r 42000_84000_M2 44000_84000_M2 0.018
r 44000_84000_M2 46000_84000_M2 0.018
r 46000_84000_M2 48000_84000_M2 0.018
r 48000_84000_M2 50000_84000_M2 0.018
r 50000_84000_M2 52000_84000_M2 0.018
r 52000_84000_M2 54000_84000_M2 0.018
r 54000_84000_M2 56000_84000_M2 0.018
r 56000_84000_M2 58000_84000_M2 0.018
r 58000_84000_M2 60000_84000_M2 0.018
r 60000_84000_M2 62000_84000_M2 0.018
r 62000_84000_M2 64000_84000_M2 0.018
r 64000_84000_M2 66000_84000_M2 0.018
r 66000_84000_M2 68000_84000_M2 0.018
r 68000_84000_M2 70000_84000_M2 0.018
r 70000_84000_M2 72000_84000_M2 0.018
r 72000_84000_M2 74000_84000_M2 0.018
r 74000_84000_M2 76000_84000_M2 0.018
r 76000_84000_M2 78000_84000_M2 0.018
r 78000_84000_M2 80000_84000_M2 0.018
r 80000_84000_M2 82000_84000_M2 0.018
r 82000_84000_M2 84000_84000_M2 0.018
r 84000_84000_M2 86000_84000_M2 0.018
r 86000_84000_M2 88000_84000_M2 0.018
r 88000_84000_M2 90000_84000_M2 0.018
r 90000_84000_M2 92000_84000_M2 0.018
r 92000_84000_M2 94000_84000_M2 0.018
r 94000_84000_M2 96000_84000_M2 0.018
r 96000_84000_M2 98000_84000_M2 0.018
r 98000_84000_M2 100000_84000_M2 0.018
r 2000_86000_M2 4000_86000_M2 0.018
r 4000_86000_M2 6000_86000_M2 0.018
r 6000_86000_M2 8000_86000_M2 0.018
r 8000_86000_M2 10000_86000_M2 0.018
r 10000_86000_M2 12000_86000_M2 0.018
r 12000_86000_M2 14000_86000_M2 0.018
r 14000_86000_M2 16000_86000_M2 0.018
r 16000_86000_M2 18000_86000_M2 0.018
r 18000_86000_M2 20000_86000_M2 0.018
r 20000_86000_M2 22000_86000_M2 0.018
r 22000_86000_M2 24000_86000_M2 0.018
r 24000_86000_M2 26000_86000_M2 0.018
r 26000_86000_M2 28000_86000_M2 0.018
r 28000_86000_M2 30000_86000_M2 0.018
r 30000_86000_M2 32000_86000_M2 0.018
r 32000_86000_M2 34000_86000_M2 0.018
r 34000_86000_M2 36000_86000_M2 0.018
r 36000_86000_M2 38000_86000_M2 0.018
r 38000_86000_M2 40000_86000_M2 0.018
r 40000_86000_M2 42000_86000_M2 0.018
r 42000_86000_M2 44000_86000_M2 0.018
r 44000_86000_M2 46000_86000_M2 0.018
r 46000_86000_M2 48000_86000_M2 0.018
r 48000_86000_M2 50000_86000_M2 0.018
r 50000_86000_M2 52000_86000_M2 0.018
r 52000_86000_M2 54000_86000_M2 0.018
r 54000_86000_M2 56000_86000_M2 0.018
r 56000_86000_M2 58000_86000_M2 0.018
r 58000_86000_M2 60000_86000_M2 0.018
r 60000_86000_M2 62000_86000_M2 0.018
r 62000_86000_M2 64000_86000_M2 0.018
r 64000_86000_M2 66000_86000_M2 0.018
r 66000_86000_M2 68000_86000_M2 0.018
r 68000_86000_M2 70000_86000_M2 0.018
r 70000_86000_M2 72000_86000_M2 0.018
r 72000_86000_M2 74000_86000_M2 0.018
r 74000_86000_M2 76000_86000_M2 0.018
r 76000_86000_M2 78000_86000_M2 0.018
r 78000_86000_M2 80000_86000_M2 0.018
r 80000_86000_M2 82000_86000_M2 0.018
r 82000_86000_M2 84000_86000_M2 0.018
r 84000_86000_M2 86000_86000_M2 0.018
r 86000_86000_M2 88000_86000_M2 0.018
r 88000_86000_M2 90000_86000_M2 0.018
r 90000_86000_M2 92000_86000_M2 0.018
r 92000_86000_M2 94000_86000_M2 0.018
r 94000_86000_M2 96000_86000_M2 0.018
r 96000_86000_M2 98000_86000_M2 0.018
r 98000_86000_M2 100000_86000_M2 0.018
r 2000_88000_M2 4000_88000_M2 0.018
r 4000_88000_M2 6000_88000_M2 0.018
r 6000_88000_M2 8000_88000_M2 0.018
r 8000_88000_M2 10000_88000_M2 0.018
r 10000_88000_M2 12000_88000_M2 0.018
r 12000_88000_M2 14000_88000_M2 0.018
r 14000_88000_M2 16000_88000_M2 0.018
r 16000_88000_M2 18000_88000_M2 0.018
r 18000_88000_M2 20000_88000_M2 0.018
r 20000_88000_M2 22000_88000_M2 0.018
r 22000_88000_M2 24000_88000_M2 0.018
r 24000_88000_M2 26000_88000_M2 0.018
r 26000_88000_M2 28000_88000_M2 0.018
r 28000_88000_M2 30000_88000_M2 0.018
r 30000_88000_M2 32000_88000_M2 0.018
r 32000_88000_M2 34000_88000_M2 0.018
r 34000_88000_M2 36000_88000_M2 0.018
r 36000_88000_M2 38000_88000_M2 0.018
r 38000_88000_M2 40000_88000_M2 0.018
r 40000_88000_M2 42000_88000_M2 0.018
r 42000_88000_M2 44000_88000_M2 0.018
r 44000_88000_M2 46000_88000_M2 0.018
r 46000_88000_M2 48000_88000_M2 0.018
r 48000_88000_M2 50000_88000_M2 0.018
r 50000_88000_M2 52000_88000_M2 0.018
r 52000_88000_M2 54000_88000_M2 0.018
r 54000_88000_M2 56000_88000_M2 0.018
r 56000_88000_M2 58000_88000_M2 0.018
r 58000_88000_M2 60000_88000_M2 0.018
r 60000_88000_M2 62000_88000_M2 0.018
r 62000_88000_M2 64000_88000_M2 0.018
r 64000_88000_M2 66000_88000_M2 0.018
r 66000_88000_M2 68000_88000_M2 0.018
r 68000_88000_M2 70000_88000_M2 0.018
r 70000_88000_M2 72000_88000_M2 0.018
r 72000_88000_M2 74000_88000_M2 0.018
r 74000_88000_M2 76000_88000_M2 0.018
r 76000_88000_M2 78000_88000_M2 0.018
r 78000_88000_M2 80000_88000_M2 0.018
r 80000_88000_M2 82000_88000_M2 0.018
r 82000_88000_M2 84000_88000_M2 0.018
r 84000_88000_M2 86000_88000_M2 0.018
r 86000_88000_M2 88000_88000_M2 0.018
r 88000_88000_M2 90000_88000_M2 0.018
r 90000_88000_M2 92000_88000_M2 0.018
r 92000_88000_M2 94000_88000_M2 0.018
r 94000_88000_M2 96000_88000_M2 0.018
r 96000_88000_M2 98000_88000_M2 0.018
r 98000_88000_M2 100000_88000_M2 0.018
r 2000_90000_M2 4000_90000_M2 0.018
r 4000_90000_M2 6000_90000_M2 0.018
r 6000_90000_M2 8000_90000_M2 0.018
r 8000_90000_M2 10000_90000_M2 0.018
r 10000_90000_M2 12000_90000_M2 0.018
r 12000_90000_M2 14000_90000_M2 0.018
r 14000_90000_M2 16000_90000_M2 0.018
r 16000_90000_M2 18000_90000_M2 0.018
r 18000_90000_M2 20000_90000_M2 0.018
r 20000_90000_M2 22000_90000_M2 0.018
r 22000_90000_M2 24000_90000_M2 0.018
r 24000_90000_M2 26000_90000_M2 0.018
r 26000_90000_M2 28000_90000_M2 0.018
r 28000_90000_M2 30000_90000_M2 0.018
r 30000_90000_M2 32000_90000_M2 0.018
r 32000_90000_M2 34000_90000_M2 0.018
r 34000_90000_M2 36000_90000_M2 0.018
r 36000_90000_M2 38000_90000_M2 0.018
r 38000_90000_M2 40000_90000_M2 0.018
r 40000_90000_M2 42000_90000_M2 0.018
r 42000_90000_M2 44000_90000_M2 0.018
r 44000_90000_M2 46000_90000_M2 0.018
r 46000_90000_M2 48000_90000_M2 0.018
r 48000_90000_M2 50000_90000_M2 0.018
r 50000_90000_M2 52000_90000_M2 0.018
r 52000_90000_M2 54000_90000_M2 0.018
r 54000_90000_M2 56000_90000_M2 0.018
r 56000_90000_M2 58000_90000_M2 0.018
r 58000_90000_M2 60000_90000_M2 0.018
r 60000_90000_M2 62000_90000_M2 0.018
r 62000_90000_M2 64000_90000_M2 0.018
r 64000_90000_M2 66000_90000_M2 0.018
r 66000_90000_M2 68000_90000_M2 0.018
r 68000_90000_M2 70000_90000_M2 0.018
r 70000_90000_M2 72000_90000_M2 0.018
r 72000_90000_M2 74000_90000_M2 0.018
r 74000_90000_M2 76000_90000_M2 0.018
r 76000_90000_M2 78000_90000_M2 0.018
r 78000_90000_M2 80000_90000_M2 0.018
r 80000_90000_M2 82000_90000_M2 0.018
r 82000_90000_M2 84000_90000_M2 0.018
r 84000_90000_M2 86000_90000_M2 0.018
r 86000_90000_M2 88000_90000_M2 0.018
r 88000_90000_M2 90000_90000_M2 0.018
r 90000_90000_M2 92000_90000_M2 0.018
r 92000_90000_M2 94000_90000_M2 0.018
r 94000_90000_M2 96000_90000_M2 0.018
r 96000_90000_M2 98000_90000_M2 0.018
r 98000_90000_M2 100000_90000_M2 0.018
r 2000_92000_M2 4000_92000_M2 0.018
r 4000_92000_M2 6000_92000_M2 0.018
r 6000_92000_M2 8000_92000_M2 0.018
r 8000_92000_M2 10000_92000_M2 0.018
r 10000_92000_M2 12000_92000_M2 0.018
r 12000_92000_M2 14000_92000_M2 0.018
r 14000_92000_M2 16000_92000_M2 0.018
r 16000_92000_M2 18000_92000_M2 0.018
r 18000_92000_M2 20000_92000_M2 0.018
r 20000_92000_M2 22000_92000_M2 0.018
r 22000_92000_M2 24000_92000_M2 0.018
r 24000_92000_M2 26000_92000_M2 0.018
r 26000_92000_M2 28000_92000_M2 0.018
r 28000_92000_M2 30000_92000_M2 0.018
r 30000_92000_M2 32000_92000_M2 0.018
r 32000_92000_M2 34000_92000_M2 0.018
r 34000_92000_M2 36000_92000_M2 0.018
r 36000_92000_M2 38000_92000_M2 0.018
r 38000_92000_M2 40000_92000_M2 0.018
r 40000_92000_M2 42000_92000_M2 0.018
r 42000_92000_M2 44000_92000_M2 0.018
r 44000_92000_M2 46000_92000_M2 0.018
r 46000_92000_M2 48000_92000_M2 0.018
r 48000_92000_M2 50000_92000_M2 0.018
r 50000_92000_M2 52000_92000_M2 0.018
r 52000_92000_M2 54000_92000_M2 0.018
r 54000_92000_M2 56000_92000_M2 0.018
r 56000_92000_M2 58000_92000_M2 0.018
r 58000_92000_M2 60000_92000_M2 0.018
r 60000_92000_M2 62000_92000_M2 0.018
r 62000_92000_M2 64000_92000_M2 0.018
r 64000_92000_M2 66000_92000_M2 0.018
r 66000_92000_M2 68000_92000_M2 0.018
r 68000_92000_M2 70000_92000_M2 0.018
r 70000_92000_M2 72000_92000_M2 0.018
r 72000_92000_M2 74000_92000_M2 0.018
r 74000_92000_M2 76000_92000_M2 0.018
r 76000_92000_M2 78000_92000_M2 0.018
r 78000_92000_M2 80000_92000_M2 0.018
r 80000_92000_M2 82000_92000_M2 0.018
r 82000_92000_M2 84000_92000_M2 0.018
r 84000_92000_M2 86000_92000_M2 0.018
r 86000_92000_M2 88000_92000_M2 0.018
r 88000_92000_M2 90000_92000_M2 0.018
r 90000_92000_M2 92000_92000_M2 0.018
r 92000_92000_M2 94000_92000_M2 0.018
r 94000_92000_M2 96000_92000_M2 0.018
r 96000_92000_M2 98000_92000_M2 0.018
r 98000_92000_M2 100000_92000_M2 0.018
r 2000_94000_M2 4000_94000_M2 0.018
r 4000_94000_M2 6000_94000_M2 0.018
r 6000_94000_M2 8000_94000_M2 0.018
r 8000_94000_M2 10000_94000_M2 0.018
r 10000_94000_M2 12000_94000_M2 0.018
r 12000_94000_M2 14000_94000_M2 0.018
r 14000_94000_M2 16000_94000_M2 0.018
r 16000_94000_M2 18000_94000_M2 0.018
r 18000_94000_M2 20000_94000_M2 0.018
r 20000_94000_M2 22000_94000_M2 0.018
r 22000_94000_M2 24000_94000_M2 0.018
r 24000_94000_M2 26000_94000_M2 0.018
r 26000_94000_M2 28000_94000_M2 0.018
r 28000_94000_M2 30000_94000_M2 0.018
r 30000_94000_M2 32000_94000_M2 0.018
r 32000_94000_M2 34000_94000_M2 0.018
r 34000_94000_M2 36000_94000_M2 0.018
r 36000_94000_M2 38000_94000_M2 0.018
r 38000_94000_M2 40000_94000_M2 0.018
r 40000_94000_M2 42000_94000_M2 0.018
r 42000_94000_M2 44000_94000_M2 0.018
r 44000_94000_M2 46000_94000_M2 0.018
r 46000_94000_M2 48000_94000_M2 0.018
r 48000_94000_M2 50000_94000_M2 0.018
r 50000_94000_M2 52000_94000_M2 0.018
r 52000_94000_M2 54000_94000_M2 0.018
r 54000_94000_M2 56000_94000_M2 0.018
r 56000_94000_M2 58000_94000_M2 0.018
r 58000_94000_M2 60000_94000_M2 0.018
r 60000_94000_M2 62000_94000_M2 0.018
r 62000_94000_M2 64000_94000_M2 0.018
r 64000_94000_M2 66000_94000_M2 0.018
r 66000_94000_M2 68000_94000_M2 0.018
r 68000_94000_M2 70000_94000_M2 0.018
r 70000_94000_M2 72000_94000_M2 0.018
r 72000_94000_M2 74000_94000_M2 0.018
r 74000_94000_M2 76000_94000_M2 0.018
r 76000_94000_M2 78000_94000_M2 0.018
r 78000_94000_M2 80000_94000_M2 0.018
r 80000_94000_M2 82000_94000_M2 0.018
r 82000_94000_M2 84000_94000_M2 0.018
r 84000_94000_M2 86000_94000_M2 0.018
r 86000_94000_M2 88000_94000_M2 0.018
r 88000_94000_M2 90000_94000_M2 0.018
r 90000_94000_M2 92000_94000_M2 0.018
r 92000_94000_M2 94000_94000_M2 0.018
r 94000_94000_M2 96000_94000_M2 0.018
r 96000_94000_M2 98000_94000_M2 0.018
r 98000_94000_M2 100000_94000_M2 0.018
r 2000_96000_M2 4000_96000_M2 0.018
r 4000_96000_M2 6000_96000_M2 0.018
r 6000_96000_M2 8000_96000_M2 0.018
r 8000_96000_M2 10000_96000_M2 0.018
r 10000_96000_M2 12000_96000_M2 0.018
r 12000_96000_M2 14000_96000_M2 0.018
r 14000_96000_M2 16000_96000_M2 0.018
r 16000_96000_M2 18000_96000_M2 0.018
r 18000_96000_M2 20000_96000_M2 0.018
r 20000_96000_M2 22000_96000_M2 0.018
r 22000_96000_M2 24000_96000_M2 0.018
r 24000_96000_M2 26000_96000_M2 0.018
r 26000_96000_M2 28000_96000_M2 0.018
r 28000_96000_M2 30000_96000_M2 0.018
r 30000_96000_M2 32000_96000_M2 0.018
r 32000_96000_M2 34000_96000_M2 0.018
r 34000_96000_M2 36000_96000_M2 0.018
r 36000_96000_M2 38000_96000_M2 0.018
r 38000_96000_M2 40000_96000_M2 0.018
r 40000_96000_M2 42000_96000_M2 0.018
r 42000_96000_M2 44000_96000_M2 0.018
r 44000_96000_M2 46000_96000_M2 0.018
r 46000_96000_M2 48000_96000_M2 0.018
r 48000_96000_M2 50000_96000_M2 0.018
r 50000_96000_M2 52000_96000_M2 0.018
r 52000_96000_M2 54000_96000_M2 0.018
r 54000_96000_M2 56000_96000_M2 0.018
r 56000_96000_M2 58000_96000_M2 0.018
r 58000_96000_M2 60000_96000_M2 0.018
r 60000_96000_M2 62000_96000_M2 0.018
r 62000_96000_M2 64000_96000_M2 0.018
r 64000_96000_M2 66000_96000_M2 0.018
r 66000_96000_M2 68000_96000_M2 0.018
r 68000_96000_M2 70000_96000_M2 0.018
r 70000_96000_M2 72000_96000_M2 0.018
r 72000_96000_M2 74000_96000_M2 0.018
r 74000_96000_M2 76000_96000_M2 0.018
r 76000_96000_M2 78000_96000_M2 0.018
r 78000_96000_M2 80000_96000_M2 0.018
r 80000_96000_M2 82000_96000_M2 0.018
r 82000_96000_M2 84000_96000_M2 0.018
r 84000_96000_M2 86000_96000_M2 0.018
r 86000_96000_M2 88000_96000_M2 0.018
r 88000_96000_M2 90000_96000_M2 0.018
r 90000_96000_M2 92000_96000_M2 0.018
r 92000_96000_M2 94000_96000_M2 0.018
r 94000_96000_M2 96000_96000_M2 0.018
r 96000_96000_M2 98000_96000_M2 0.018
r 98000_96000_M2 100000_96000_M2 0.018
r 2000_98000_M2 4000_98000_M2 0.018
r 4000_98000_M2 6000_98000_M2 0.018
r 6000_98000_M2 8000_98000_M2 0.018
r 8000_98000_M2 10000_98000_M2 0.018
r 10000_98000_M2 12000_98000_M2 0.018
r 12000_98000_M2 14000_98000_M2 0.018
r 14000_98000_M2 16000_98000_M2 0.018
r 16000_98000_M2 18000_98000_M2 0.018
r 18000_98000_M2 20000_98000_M2 0.018
r 20000_98000_M2 22000_98000_M2 0.018
r 22000_98000_M2 24000_98000_M2 0.018
r 24000_98000_M2 26000_98000_M2 0.018
r 26000_98000_M2 28000_98000_M2 0.018
r 28000_98000_M2 30000_98000_M2 0.018
r 30000_98000_M2 32000_98000_M2 0.018
r 32000_98000_M2 34000_98000_M2 0.018
r 34000_98000_M2 36000_98000_M2 0.018
r 36000_98000_M2 38000_98000_M2 0.018
r 38000_98000_M2 40000_98000_M2 0.018
r 40000_98000_M2 42000_98000_M2 0.018
r 42000_98000_M2 44000_98000_M2 0.018
r 44000_98000_M2 46000_98000_M2 0.018
r 46000_98000_M2 48000_98000_M2 0.018
r 48000_98000_M2 50000_98000_M2 0.018
r 50000_98000_M2 52000_98000_M2 0.018
r 52000_98000_M2 54000_98000_M2 0.018
r 54000_98000_M2 56000_98000_M2 0.018
r 56000_98000_M2 58000_98000_M2 0.018
r 58000_98000_M2 60000_98000_M2 0.018
r 60000_98000_M2 62000_98000_M2 0.018
r 62000_98000_M2 64000_98000_M2 0.018
r 64000_98000_M2 66000_98000_M2 0.018
r 66000_98000_M2 68000_98000_M2 0.018
r 68000_98000_M2 70000_98000_M2 0.018
r 70000_98000_M2 72000_98000_M2 0.018
r 72000_98000_M2 74000_98000_M2 0.018
r 74000_98000_M2 76000_98000_M2 0.018
r 76000_98000_M2 78000_98000_M2 0.018
r 78000_98000_M2 80000_98000_M2 0.018
r 80000_98000_M2 82000_98000_M2 0.018
r 82000_98000_M2 84000_98000_M2 0.018
r 84000_98000_M2 86000_98000_M2 0.018
r 86000_98000_M2 88000_98000_M2 0.018
r 88000_98000_M2 90000_98000_M2 0.018
r 90000_98000_M2 92000_98000_M2 0.018
r 92000_98000_M2 94000_98000_M2 0.018
r 94000_98000_M2 96000_98000_M2 0.018
r 96000_98000_M2 98000_98000_M2 0.018
r 98000_98000_M2 100000_98000_M2 0.018
r 2000_100000_M2 4000_100000_M2 0.018
r 4000_100000_M2 6000_100000_M2 0.018
r 6000_100000_M2 8000_100000_M2 0.018
r 8000_100000_M2 10000_100000_M2 0.018
r 10000_100000_M2 12000_100000_M2 0.018
r 12000_100000_M2 14000_100000_M2 0.018
r 14000_100000_M2 16000_100000_M2 0.018
r 16000_100000_M2 18000_100000_M2 0.018
r 18000_100000_M2 20000_100000_M2 0.018
r 20000_100000_M2 22000_100000_M2 0.018
r 22000_100000_M2 24000_100000_M2 0.018
r 24000_100000_M2 26000_100000_M2 0.018
r 26000_100000_M2 28000_100000_M2 0.018
r 28000_100000_M2 30000_100000_M2 0.018
r 30000_100000_M2 32000_100000_M2 0.018
r 32000_100000_M2 34000_100000_M2 0.018
r 34000_100000_M2 36000_100000_M2 0.018
r 36000_100000_M2 38000_100000_M2 0.018
r 38000_100000_M2 40000_100000_M2 0.018
r 40000_100000_M2 42000_100000_M2 0.018
r 42000_100000_M2 44000_100000_M2 0.018
r 44000_100000_M2 46000_100000_M2 0.018
r 46000_100000_M2 48000_100000_M2 0.018
r 48000_100000_M2 50000_100000_M2 0.018
r 50000_100000_M2 52000_100000_M2 0.018
r 52000_100000_M2 54000_100000_M2 0.018
r 54000_100000_M2 56000_100000_M2 0.018
r 56000_100000_M2 58000_100000_M2 0.018
r 58000_100000_M2 60000_100000_M2 0.018
r 60000_100000_M2 62000_100000_M2 0.018
r 62000_100000_M2 64000_100000_M2 0.018
r 64000_100000_M2 66000_100000_M2 0.018
r 66000_100000_M2 68000_100000_M2 0.018
r 68000_100000_M2 70000_100000_M2 0.018
r 70000_100000_M2 72000_100000_M2 0.018
r 72000_100000_M2 74000_100000_M2 0.018
r 74000_100000_M2 76000_100000_M2 0.018
r 76000_100000_M2 78000_100000_M2 0.018
r 78000_100000_M2 80000_100000_M2 0.018
r 80000_100000_M2 82000_100000_M2 0.018
r 82000_100000_M2 84000_100000_M2 0.018
r 84000_100000_M2 86000_100000_M2 0.018
r 86000_100000_M2 88000_100000_M2 0.018
r 88000_100000_M2 90000_100000_M2 0.018
r 90000_100000_M2 92000_100000_M2 0.018
r 92000_100000_M2 94000_100000_M2 0.018
r 94000_100000_M2 96000_100000_M2 0.018
r 96000_100000_M2 98000_100000_M2 0.018
r 98000_100000_M2 100000_100000_M2 0.018

* M2 Vertical resistors
r 2000_2000_M2 2000_4000_M2 0.022
r 2000_4000_M2 2000_6000_M2 0.022
r 2000_6000_M2 2000_8000_M2 0.022
r 2000_8000_M2 2000_10000_M2 0.022
r 2000_10000_M2 2000_12000_M2 0.022
r 2000_12000_M2 2000_14000_M2 0.022
r 2000_14000_M2 2000_16000_M2 0.022
r 2000_16000_M2 2000_18000_M2 0.022
r 2000_18000_M2 2000_20000_M2 0.022
r 2000_20000_M2 2000_22000_M2 0.022
r 2000_22000_M2 2000_24000_M2 0.022
r 2000_24000_M2 2000_26000_M2 0.022
r 2000_26000_M2 2000_28000_M2 0.022
r 2000_28000_M2 2000_30000_M2 0.022
r 2000_30000_M2 2000_32000_M2 0.022
r 2000_32000_M2 2000_34000_M2 0.022
r 2000_34000_M2 2000_36000_M2 0.022
r 2000_36000_M2 2000_38000_M2 0.022
r 2000_38000_M2 2000_40000_M2 0.022
r 2000_40000_M2 2000_42000_M2 0.022
r 2000_42000_M2 2000_44000_M2 0.022
r 2000_44000_M2 2000_46000_M2 0.022
r 2000_46000_M2 2000_48000_M2 0.022
r 2000_48000_M2 2000_50000_M2 0.022
r 2000_50000_M2 2000_52000_M2 0.022
r 2000_52000_M2 2000_54000_M2 0.022
r 2000_54000_M2 2000_56000_M2 0.022
r 2000_56000_M2 2000_58000_M2 0.022
r 2000_58000_M2 2000_60000_M2 0.022
r 2000_60000_M2 2000_62000_M2 0.022
r 2000_62000_M2 2000_64000_M2 0.022
r 2000_64000_M2 2000_66000_M2 0.022
r 2000_66000_M2 2000_68000_M2 0.022
r 2000_68000_M2 2000_70000_M2 0.022
r 2000_70000_M2 2000_72000_M2 0.022
r 2000_72000_M2 2000_74000_M2 0.022
r 2000_74000_M2 2000_76000_M2 0.022
r 2000_76000_M2 2000_78000_M2 0.022
r 2000_78000_M2 2000_80000_M2 0.022
r 2000_80000_M2 2000_82000_M2 0.022
r 2000_82000_M2 2000_84000_M2 0.022
r 2000_84000_M2 2000_86000_M2 0.022
r 2000_86000_M2 2000_88000_M2 0.022
r 2000_88000_M2 2000_90000_M2 0.022
r 2000_90000_M2 2000_92000_M2 0.022
r 2000_92000_M2 2000_94000_M2 0.022
r 2000_94000_M2 2000_96000_M2 0.022
r 2000_96000_M2 2000_98000_M2 0.022
r 2000_98000_M2 2000_100000_M2 0.022
r 4000_2000_M2 4000_4000_M2 0.022
r 4000_4000_M2 4000_6000_M2 0.022
r 4000_6000_M2 4000_8000_M2 0.022
r 4000_8000_M2 4000_10000_M2 0.022
r 4000_10000_M2 4000_12000_M2 0.022
r 4000_12000_M2 4000_14000_M2 0.022
r 4000_14000_M2 4000_16000_M2 0.022
r 4000_16000_M2 4000_18000_M2 0.022
r 4000_18000_M2 4000_20000_M2 0.022
r 4000_20000_M2 4000_22000_M2 0.022
r 4000_22000_M2 4000_24000_M2 0.022
r 4000_24000_M2 4000_26000_M2 0.022
r 4000_26000_M2 4000_28000_M2 0.022
r 4000_28000_M2 4000_30000_M2 0.022
r 4000_30000_M2 4000_32000_M2 0.022
r 4000_32000_M2 4000_34000_M2 0.022
r 4000_34000_M2 4000_36000_M2 0.022
r 4000_36000_M2 4000_38000_M2 0.022
r 4000_38000_M2 4000_40000_M2 0.022
r 4000_40000_M2 4000_42000_M2 0.022
r 4000_42000_M2 4000_44000_M2 0.022
r 4000_44000_M2 4000_46000_M2 0.022
r 4000_46000_M2 4000_48000_M2 0.022
r 4000_48000_M2 4000_50000_M2 0.022
r 4000_50000_M2 4000_52000_M2 0.022
r 4000_52000_M2 4000_54000_M2 0.022
r 4000_54000_M2 4000_56000_M2 0.022
r 4000_56000_M2 4000_58000_M2 0.022
r 4000_58000_M2 4000_60000_M2 0.022
r 4000_60000_M2 4000_62000_M2 0.022
r 4000_62000_M2 4000_64000_M2 0.022
r 4000_64000_M2 4000_66000_M2 0.022
r 4000_66000_M2 4000_68000_M2 0.022
r 4000_68000_M2 4000_70000_M2 0.022
r 4000_70000_M2 4000_72000_M2 0.022
r 4000_72000_M2 4000_74000_M2 0.022
r 4000_74000_M2 4000_76000_M2 0.022
r 4000_76000_M2 4000_78000_M2 0.022
r 4000_78000_M2 4000_80000_M2 0.022
r 4000_80000_M2 4000_82000_M2 0.022
r 4000_82000_M2 4000_84000_M2 0.022
r 4000_84000_M2 4000_86000_M2 0.022
r 4000_86000_M2 4000_88000_M2 0.022
r 4000_88000_M2 4000_90000_M2 0.022
r 4000_90000_M2 4000_92000_M2 0.022
r 4000_92000_M2 4000_94000_M2 0.022
r 4000_94000_M2 4000_96000_M2 0.022
r 4000_96000_M2 4000_98000_M2 0.022
r 4000_98000_M2 4000_100000_M2 0.022
r 6000_2000_M2 6000_4000_M2 0.022
r 6000_4000_M2 6000_6000_M2 0.022
r 6000_6000_M2 6000_8000_M2 0.022
r 6000_8000_M2 6000_10000_M2 0.022
r 6000_10000_M2 6000_12000_M2 0.022
r 6000_12000_M2 6000_14000_M2 0.022
r 6000_14000_M2 6000_16000_M2 0.022
r 6000_16000_M2 6000_18000_M2 0.022
r 6000_18000_M2 6000_20000_M2 0.022
r 6000_20000_M2 6000_22000_M2 0.022
r 6000_22000_M2 6000_24000_M2 0.022
r 6000_24000_M2 6000_26000_M2 0.022
r 6000_26000_M2 6000_28000_M2 0.022
r 6000_28000_M2 6000_30000_M2 0.022
r 6000_30000_M2 6000_32000_M2 0.022
r 6000_32000_M2 6000_34000_M2 0.022
r 6000_34000_M2 6000_36000_M2 0.022
r 6000_36000_M2 6000_38000_M2 0.022
r 6000_38000_M2 6000_40000_M2 0.022
r 6000_40000_M2 6000_42000_M2 0.022
r 6000_42000_M2 6000_44000_M2 0.022
r 6000_44000_M2 6000_46000_M2 0.022
r 6000_46000_M2 6000_48000_M2 0.022
r 6000_48000_M2 6000_50000_M2 0.022
r 6000_50000_M2 6000_52000_M2 0.022
r 6000_52000_M2 6000_54000_M2 0.022
r 6000_54000_M2 6000_56000_M2 0.022
r 6000_56000_M2 6000_58000_M2 0.022
r 6000_58000_M2 6000_60000_M2 0.022
r 6000_60000_M2 6000_62000_M2 0.022
r 6000_62000_M2 6000_64000_M2 0.022
r 6000_64000_M2 6000_66000_M2 0.022
r 6000_66000_M2 6000_68000_M2 0.022
r 6000_68000_M2 6000_70000_M2 0.022
r 6000_70000_M2 6000_72000_M2 0.022
r 6000_72000_M2 6000_74000_M2 0.022
r 6000_74000_M2 6000_76000_M2 0.022
r 6000_76000_M2 6000_78000_M2 0.022
r 6000_78000_M2 6000_80000_M2 0.022
r 6000_80000_M2 6000_82000_M2 0.022
r 6000_82000_M2 6000_84000_M2 0.022
r 6000_84000_M2 6000_86000_M2 0.022
r 6000_86000_M2 6000_88000_M2 0.022
r 6000_88000_M2 6000_90000_M2 0.022
r 6000_90000_M2 6000_92000_M2 0.022
r 6000_92000_M2 6000_94000_M2 0.022
r 6000_94000_M2 6000_96000_M2 0.022
r 6000_96000_M2 6000_98000_M2 0.022
r 6000_98000_M2 6000_100000_M2 0.022
r 8000_2000_M2 8000_4000_M2 0.022
r 8000_4000_M2 8000_6000_M2 0.022
r 8000_6000_M2 8000_8000_M2 0.022
r 8000_8000_M2 8000_10000_M2 0.022
r 8000_10000_M2 8000_12000_M2 0.022
r 8000_12000_M2 8000_14000_M2 0.022
r 8000_14000_M2 8000_16000_M2 0.022
r 8000_16000_M2 8000_18000_M2 0.022
r 8000_18000_M2 8000_20000_M2 0.022
r 8000_20000_M2 8000_22000_M2 0.022
r 8000_22000_M2 8000_24000_M2 0.022
r 8000_24000_M2 8000_26000_M2 0.022
r 8000_26000_M2 8000_28000_M2 0.022
r 8000_28000_M2 8000_30000_M2 0.022
r 8000_30000_M2 8000_32000_M2 0.022
r 8000_32000_M2 8000_34000_M2 0.022
r 8000_34000_M2 8000_36000_M2 0.022
r 8000_36000_M2 8000_38000_M2 0.022
r 8000_38000_M2 8000_40000_M2 0.022
r 8000_40000_M2 8000_42000_M2 0.022
r 8000_42000_M2 8000_44000_M2 0.022
r 8000_44000_M2 8000_46000_M2 0.022
r 8000_46000_M2 8000_48000_M2 0.022
r 8000_48000_M2 8000_50000_M2 0.022
r 8000_50000_M2 8000_52000_M2 0.022
r 8000_52000_M2 8000_54000_M2 0.022
r 8000_54000_M2 8000_56000_M2 0.022
r 8000_56000_M2 8000_58000_M2 0.022
r 8000_58000_M2 8000_60000_M2 0.022
r 8000_60000_M2 8000_62000_M2 0.022
r 8000_62000_M2 8000_64000_M2 0.022
r 8000_64000_M2 8000_66000_M2 0.022
r 8000_66000_M2 8000_68000_M2 0.022
r 8000_68000_M2 8000_70000_M2 0.022
r 8000_70000_M2 8000_72000_M2 0.022
r 8000_72000_M2 8000_74000_M2 0.022
r 8000_74000_M2 8000_76000_M2 0.022
r 8000_76000_M2 8000_78000_M2 0.022
r 8000_78000_M2 8000_80000_M2 0.022
r 8000_80000_M2 8000_82000_M2 0.022
r 8000_82000_M2 8000_84000_M2 0.022
r 8000_84000_M2 8000_86000_M2 0.022
r 8000_86000_M2 8000_88000_M2 0.022
r 8000_88000_M2 8000_90000_M2 0.022
r 8000_90000_M2 8000_92000_M2 0.022
r 8000_92000_M2 8000_94000_M2 0.022
r 8000_94000_M2 8000_96000_M2 0.022
r 8000_96000_M2 8000_98000_M2 0.022
r 8000_98000_M2 8000_100000_M2 0.022
r 10000_2000_M2 10000_4000_M2 0.022
r 10000_4000_M2 10000_6000_M2 0.022
r 10000_6000_M2 10000_8000_M2 0.022
r 10000_8000_M2 10000_10000_M2 0.022
r 10000_10000_M2 10000_12000_M2 0.022
r 10000_12000_M2 10000_14000_M2 0.022
r 10000_14000_M2 10000_16000_M2 0.022
r 10000_16000_M2 10000_18000_M2 0.022
r 10000_18000_M2 10000_20000_M2 0.022
r 10000_20000_M2 10000_22000_M2 0.022
r 10000_22000_M2 10000_24000_M2 0.022
r 10000_24000_M2 10000_26000_M2 0.022
r 10000_26000_M2 10000_28000_M2 0.022
r 10000_28000_M2 10000_30000_M2 0.022
r 10000_30000_M2 10000_32000_M2 0.022
r 10000_32000_M2 10000_34000_M2 0.022
r 10000_34000_M2 10000_36000_M2 0.022
r 10000_36000_M2 10000_38000_M2 0.022
r 10000_38000_M2 10000_40000_M2 0.022
r 10000_40000_M2 10000_42000_M2 0.022
r 10000_42000_M2 10000_44000_M2 0.022
r 10000_44000_M2 10000_46000_M2 0.022
r 10000_46000_M2 10000_48000_M2 0.022
r 10000_48000_M2 10000_50000_M2 0.022
r 10000_50000_M2 10000_52000_M2 0.022
r 10000_52000_M2 10000_54000_M2 0.022
r 10000_54000_M2 10000_56000_M2 0.022
r 10000_56000_M2 10000_58000_M2 0.022
r 10000_58000_M2 10000_60000_M2 0.022
r 10000_60000_M2 10000_62000_M2 0.022
r 10000_62000_M2 10000_64000_M2 0.022
r 10000_64000_M2 10000_66000_M2 0.022
r 10000_66000_M2 10000_68000_M2 0.022
r 10000_68000_M2 10000_70000_M2 0.022
r 10000_70000_M2 10000_72000_M2 0.022
r 10000_72000_M2 10000_74000_M2 0.022
r 10000_74000_M2 10000_76000_M2 0.022
r 10000_76000_M2 10000_78000_M2 0.022
r 10000_78000_M2 10000_80000_M2 0.022
r 10000_80000_M2 10000_82000_M2 0.022
r 10000_82000_M2 10000_84000_M2 0.022
r 10000_84000_M2 10000_86000_M2 0.022
r 10000_86000_M2 10000_88000_M2 0.022
r 10000_88000_M2 10000_90000_M2 0.022
r 10000_90000_M2 10000_92000_M2 0.022
r 10000_92000_M2 10000_94000_M2 0.022
r 10000_94000_M2 10000_96000_M2 0.022
r 10000_96000_M2 10000_98000_M2 0.022
r 10000_98000_M2 10000_100000_M2 0.022
r 12000_2000_M2 12000_4000_M2 0.022
r 12000_4000_M2 12000_6000_M2 0.022
r 12000_6000_M2 12000_8000_M2 0.022
r 12000_8000_M2 12000_10000_M2 0.022
r 12000_10000_M2 12000_12000_M2 0.022
r 12000_12000_M2 12000_14000_M2 0.022
r 12000_14000_M2 12000_16000_M2 0.022
r 12000_16000_M2 12000_18000_M2 0.022
r 12000_18000_M2 12000_20000_M2 0.022
r 12000_20000_M2 12000_22000_M2 0.022
r 12000_22000_M2 12000_24000_M2 0.022
r 12000_24000_M2 12000_26000_M2 0.022
r 12000_26000_M2 12000_28000_M2 0.022
r 12000_28000_M2 12000_30000_M2 0.022
r 12000_30000_M2 12000_32000_M2 0.022
r 12000_32000_M2 12000_34000_M2 0.022
r 12000_34000_M2 12000_36000_M2 0.022
r 12000_36000_M2 12000_38000_M2 0.022
r 12000_38000_M2 12000_40000_M2 0.022
r 12000_40000_M2 12000_42000_M2 0.022
r 12000_42000_M2 12000_44000_M2 0.022
r 12000_44000_M2 12000_46000_M2 0.022
r 12000_46000_M2 12000_48000_M2 0.022
r 12000_48000_M2 12000_50000_M2 0.022
r 12000_50000_M2 12000_52000_M2 0.022
r 12000_52000_M2 12000_54000_M2 0.022
r 12000_54000_M2 12000_56000_M2 0.022
r 12000_56000_M2 12000_58000_M2 0.022
r 12000_58000_M2 12000_60000_M2 0.022
r 12000_60000_M2 12000_62000_M2 0.022
r 12000_62000_M2 12000_64000_M2 0.022
r 12000_64000_M2 12000_66000_M2 0.022
r 12000_66000_M2 12000_68000_M2 0.022
r 12000_68000_M2 12000_70000_M2 0.022
r 12000_70000_M2 12000_72000_M2 0.022
r 12000_72000_M2 12000_74000_M2 0.022
r 12000_74000_M2 12000_76000_M2 0.022
r 12000_76000_M2 12000_78000_M2 0.022
r 12000_78000_M2 12000_80000_M2 0.022
r 12000_80000_M2 12000_82000_M2 0.022
r 12000_82000_M2 12000_84000_M2 0.022
r 12000_84000_M2 12000_86000_M2 0.022
r 12000_86000_M2 12000_88000_M2 0.022
r 12000_88000_M2 12000_90000_M2 0.022
r 12000_90000_M2 12000_92000_M2 0.022
r 12000_92000_M2 12000_94000_M2 0.022
r 12000_94000_M2 12000_96000_M2 0.022
r 12000_96000_M2 12000_98000_M2 0.022
r 12000_98000_M2 12000_100000_M2 0.022
r 14000_2000_M2 14000_4000_M2 0.022
r 14000_4000_M2 14000_6000_M2 0.022
r 14000_6000_M2 14000_8000_M2 0.022
r 14000_8000_M2 14000_10000_M2 0.022
r 14000_10000_M2 14000_12000_M2 0.022
r 14000_12000_M2 14000_14000_M2 0.022
r 14000_14000_M2 14000_16000_M2 0.022
r 14000_16000_M2 14000_18000_M2 0.022
r 14000_18000_M2 14000_20000_M2 0.022
r 14000_20000_M2 14000_22000_M2 0.022
r 14000_22000_M2 14000_24000_M2 0.022
r 14000_24000_M2 14000_26000_M2 0.022
r 14000_26000_M2 14000_28000_M2 0.022
r 14000_28000_M2 14000_30000_M2 0.022
r 14000_30000_M2 14000_32000_M2 0.022
r 14000_32000_M2 14000_34000_M2 0.022
r 14000_34000_M2 14000_36000_M2 0.022
r 14000_36000_M2 14000_38000_M2 0.022
r 14000_38000_M2 14000_40000_M2 0.022
r 14000_40000_M2 14000_42000_M2 0.022
r 14000_42000_M2 14000_44000_M2 0.022
r 14000_44000_M2 14000_46000_M2 0.022
r 14000_46000_M2 14000_48000_M2 0.022
r 14000_48000_M2 14000_50000_M2 0.022
r 14000_50000_M2 14000_52000_M2 0.022
r 14000_52000_M2 14000_54000_M2 0.022
r 14000_54000_M2 14000_56000_M2 0.022
r 14000_56000_M2 14000_58000_M2 0.022
r 14000_58000_M2 14000_60000_M2 0.022
r 14000_60000_M2 14000_62000_M2 0.022
r 14000_62000_M2 14000_64000_M2 0.022
r 14000_64000_M2 14000_66000_M2 0.022
r 14000_66000_M2 14000_68000_M2 0.022
r 14000_68000_M2 14000_70000_M2 0.022
r 14000_70000_M2 14000_72000_M2 0.022
r 14000_72000_M2 14000_74000_M2 0.022
r 14000_74000_M2 14000_76000_M2 0.022
r 14000_76000_M2 14000_78000_M2 0.022
r 14000_78000_M2 14000_80000_M2 0.022
r 14000_80000_M2 14000_82000_M2 0.022
r 14000_82000_M2 14000_84000_M2 0.022
r 14000_84000_M2 14000_86000_M2 0.022
r 14000_86000_M2 14000_88000_M2 0.022
r 14000_88000_M2 14000_90000_M2 0.022
r 14000_90000_M2 14000_92000_M2 0.022
r 14000_92000_M2 14000_94000_M2 0.022
r 14000_94000_M2 14000_96000_M2 0.022
r 14000_96000_M2 14000_98000_M2 0.022
r 14000_98000_M2 14000_100000_M2 0.022
r 16000_2000_M2 16000_4000_M2 0.022
r 16000_4000_M2 16000_6000_M2 0.022
r 16000_6000_M2 16000_8000_M2 0.022
r 16000_8000_M2 16000_10000_M2 0.022
r 16000_10000_M2 16000_12000_M2 0.022
r 16000_12000_M2 16000_14000_M2 0.022
r 16000_14000_M2 16000_16000_M2 0.022
r 16000_16000_M2 16000_18000_M2 0.022
r 16000_18000_M2 16000_20000_M2 0.022
r 16000_20000_M2 16000_22000_M2 0.022
r 16000_22000_M2 16000_24000_M2 0.022
r 16000_24000_M2 16000_26000_M2 0.022
r 16000_26000_M2 16000_28000_M2 0.022
r 16000_28000_M2 16000_30000_M2 0.022
r 16000_30000_M2 16000_32000_M2 0.022
r 16000_32000_M2 16000_34000_M2 0.022
r 16000_34000_M2 16000_36000_M2 0.022
r 16000_36000_M2 16000_38000_M2 0.022
r 16000_38000_M2 16000_40000_M2 0.022
r 16000_40000_M2 16000_42000_M2 0.022
r 16000_42000_M2 16000_44000_M2 0.022
r 16000_44000_M2 16000_46000_M2 0.022
r 16000_46000_M2 16000_48000_M2 0.022
r 16000_48000_M2 16000_50000_M2 0.022
r 16000_50000_M2 16000_52000_M2 0.022
r 16000_52000_M2 16000_54000_M2 0.022
r 16000_54000_M2 16000_56000_M2 0.022
r 16000_56000_M2 16000_58000_M2 0.022
r 16000_58000_M2 16000_60000_M2 0.022
r 16000_60000_M2 16000_62000_M2 0.022
r 16000_62000_M2 16000_64000_M2 0.022
r 16000_64000_M2 16000_66000_M2 0.022
r 16000_66000_M2 16000_68000_M2 0.022
r 16000_68000_M2 16000_70000_M2 0.022
r 16000_70000_M2 16000_72000_M2 0.022
r 16000_72000_M2 16000_74000_M2 0.022
r 16000_74000_M2 16000_76000_M2 0.022
r 16000_76000_M2 16000_78000_M2 0.022
r 16000_78000_M2 16000_80000_M2 0.022
r 16000_80000_M2 16000_82000_M2 0.022
r 16000_82000_M2 16000_84000_M2 0.022
r 16000_84000_M2 16000_86000_M2 0.022
r 16000_86000_M2 16000_88000_M2 0.022
r 16000_88000_M2 16000_90000_M2 0.022
r 16000_90000_M2 16000_92000_M2 0.022
r 16000_92000_M2 16000_94000_M2 0.022
r 16000_94000_M2 16000_96000_M2 0.022
r 16000_96000_M2 16000_98000_M2 0.022
r 16000_98000_M2 16000_100000_M2 0.022
r 18000_2000_M2 18000_4000_M2 0.022
r 18000_4000_M2 18000_6000_M2 0.022
r 18000_6000_M2 18000_8000_M2 0.022
r 18000_8000_M2 18000_10000_M2 0.022
r 18000_10000_M2 18000_12000_M2 0.022
r 18000_12000_M2 18000_14000_M2 0.022
r 18000_14000_M2 18000_16000_M2 0.022
r 18000_16000_M2 18000_18000_M2 0.022
r 18000_18000_M2 18000_20000_M2 0.022
r 18000_20000_M2 18000_22000_M2 0.022
r 18000_22000_M2 18000_24000_M2 0.022
r 18000_24000_M2 18000_26000_M2 0.022
r 18000_26000_M2 18000_28000_M2 0.022
r 18000_28000_M2 18000_30000_M2 0.022
r 18000_30000_M2 18000_32000_M2 0.022
r 18000_32000_M2 18000_34000_M2 0.022
r 18000_34000_M2 18000_36000_M2 0.022
r 18000_36000_M2 18000_38000_M2 0.022
r 18000_38000_M2 18000_40000_M2 0.022
r 18000_40000_M2 18000_42000_M2 0.022
r 18000_42000_M2 18000_44000_M2 0.022
r 18000_44000_M2 18000_46000_M2 0.022
r 18000_46000_M2 18000_48000_M2 0.022
r 18000_48000_M2 18000_50000_M2 0.022
r 18000_50000_M2 18000_52000_M2 0.022
r 18000_52000_M2 18000_54000_M2 0.022
r 18000_54000_M2 18000_56000_M2 0.022
r 18000_56000_M2 18000_58000_M2 0.022
r 18000_58000_M2 18000_60000_M2 0.022
r 18000_60000_M2 18000_62000_M2 0.022
r 18000_62000_M2 18000_64000_M2 0.022
r 18000_64000_M2 18000_66000_M2 0.022
r 18000_66000_M2 18000_68000_M2 0.022
r 18000_68000_M2 18000_70000_M2 0.022
r 18000_70000_M2 18000_72000_M2 0.022
r 18000_72000_M2 18000_74000_M2 0.022
r 18000_74000_M2 18000_76000_M2 0.022
r 18000_76000_M2 18000_78000_M2 0.022
r 18000_78000_M2 18000_80000_M2 0.022
r 18000_80000_M2 18000_82000_M2 0.022
r 18000_82000_M2 18000_84000_M2 0.022
r 18000_84000_M2 18000_86000_M2 0.022
r 18000_86000_M2 18000_88000_M2 0.022
r 18000_88000_M2 18000_90000_M2 0.022
r 18000_90000_M2 18000_92000_M2 0.022
r 18000_92000_M2 18000_94000_M2 0.022
r 18000_94000_M2 18000_96000_M2 0.022
r 18000_96000_M2 18000_98000_M2 0.022
r 18000_98000_M2 18000_100000_M2 0.022
r 20000_2000_M2 20000_4000_M2 0.022
r 20000_4000_M2 20000_6000_M2 0.022
r 20000_6000_M2 20000_8000_M2 0.022
r 20000_8000_M2 20000_10000_M2 0.022
r 20000_10000_M2 20000_12000_M2 0.022
r 20000_12000_M2 20000_14000_M2 0.022
r 20000_14000_M2 20000_16000_M2 0.022
r 20000_16000_M2 20000_18000_M2 0.022
r 20000_18000_M2 20000_20000_M2 0.022
r 20000_20000_M2 20000_22000_M2 0.022
r 20000_22000_M2 20000_24000_M2 0.022
r 20000_24000_M2 20000_26000_M2 0.022
r 20000_26000_M2 20000_28000_M2 0.022
r 20000_28000_M2 20000_30000_M2 0.022
r 20000_30000_M2 20000_32000_M2 0.022
r 20000_32000_M2 20000_34000_M2 0.022
r 20000_34000_M2 20000_36000_M2 0.022
r 20000_36000_M2 20000_38000_M2 0.022
r 20000_38000_M2 20000_40000_M2 0.022
r 20000_40000_M2 20000_42000_M2 0.022
r 20000_42000_M2 20000_44000_M2 0.022
r 20000_44000_M2 20000_46000_M2 0.022
r 20000_46000_M2 20000_48000_M2 0.022
r 20000_48000_M2 20000_50000_M2 0.022
r 20000_50000_M2 20000_52000_M2 0.022
r 20000_52000_M2 20000_54000_M2 0.022
r 20000_54000_M2 20000_56000_M2 0.022
r 20000_56000_M2 20000_58000_M2 0.022
r 20000_58000_M2 20000_60000_M2 0.022
r 20000_60000_M2 20000_62000_M2 0.022
r 20000_62000_M2 20000_64000_M2 0.022
r 20000_64000_M2 20000_66000_M2 0.022
r 20000_66000_M2 20000_68000_M2 0.022
r 20000_68000_M2 20000_70000_M2 0.022
r 20000_70000_M2 20000_72000_M2 0.022
r 20000_72000_M2 20000_74000_M2 0.022
r 20000_74000_M2 20000_76000_M2 0.022
r 20000_76000_M2 20000_78000_M2 0.022
r 20000_78000_M2 20000_80000_M2 0.022
r 20000_80000_M2 20000_82000_M2 0.022
r 20000_82000_M2 20000_84000_M2 0.022
r 20000_84000_M2 20000_86000_M2 0.022
r 20000_86000_M2 20000_88000_M2 0.022
r 20000_88000_M2 20000_90000_M2 0.022
r 20000_90000_M2 20000_92000_M2 0.022
r 20000_92000_M2 20000_94000_M2 0.022
r 20000_94000_M2 20000_96000_M2 0.022
r 20000_96000_M2 20000_98000_M2 0.022
r 20000_98000_M2 20000_100000_M2 0.022
r 22000_2000_M2 22000_4000_M2 0.022
r 22000_4000_M2 22000_6000_M2 0.022
r 22000_6000_M2 22000_8000_M2 0.022
r 22000_8000_M2 22000_10000_M2 0.022
r 22000_10000_M2 22000_12000_M2 0.022
r 22000_12000_M2 22000_14000_M2 0.022
r 22000_14000_M2 22000_16000_M2 0.022
r 22000_16000_M2 22000_18000_M2 0.022
r 22000_18000_M2 22000_20000_M2 0.022
r 22000_20000_M2 22000_22000_M2 0.022
r 22000_22000_M2 22000_24000_M2 0.022
r 22000_24000_M2 22000_26000_M2 0.022
r 22000_26000_M2 22000_28000_M2 0.022
r 22000_28000_M2 22000_30000_M2 0.022
r 22000_30000_M2 22000_32000_M2 0.022
r 22000_32000_M2 22000_34000_M2 0.022
r 22000_34000_M2 22000_36000_M2 0.022
r 22000_36000_M2 22000_38000_M2 0.022
r 22000_38000_M2 22000_40000_M2 0.022
r 22000_40000_M2 22000_42000_M2 0.022
r 22000_42000_M2 22000_44000_M2 0.022
r 22000_44000_M2 22000_46000_M2 0.022
r 22000_46000_M2 22000_48000_M2 0.022
r 22000_48000_M2 22000_50000_M2 0.022
r 22000_50000_M2 22000_52000_M2 0.022
r 22000_52000_M2 22000_54000_M2 0.022
r 22000_54000_M2 22000_56000_M2 0.022
r 22000_56000_M2 22000_58000_M2 0.022
r 22000_58000_M2 22000_60000_M2 0.022
r 22000_60000_M2 22000_62000_M2 0.022
r 22000_62000_M2 22000_64000_M2 0.022
r 22000_64000_M2 22000_66000_M2 0.022
r 22000_66000_M2 22000_68000_M2 0.022
r 22000_68000_M2 22000_70000_M2 0.022
r 22000_70000_M2 22000_72000_M2 0.022
r 22000_72000_M2 22000_74000_M2 0.022
r 22000_74000_M2 22000_76000_M2 0.022
r 22000_76000_M2 22000_78000_M2 0.022
r 22000_78000_M2 22000_80000_M2 0.022
r 22000_80000_M2 22000_82000_M2 0.022
r 22000_82000_M2 22000_84000_M2 0.022
r 22000_84000_M2 22000_86000_M2 0.022
r 22000_86000_M2 22000_88000_M2 0.022
r 22000_88000_M2 22000_90000_M2 0.022
r 22000_90000_M2 22000_92000_M2 0.022
r 22000_92000_M2 22000_94000_M2 0.022
r 22000_94000_M2 22000_96000_M2 0.022
r 22000_96000_M2 22000_98000_M2 0.022
r 22000_98000_M2 22000_100000_M2 0.022
r 24000_2000_M2 24000_4000_M2 0.022
r 24000_4000_M2 24000_6000_M2 0.022
r 24000_6000_M2 24000_8000_M2 0.022
r 24000_8000_M2 24000_10000_M2 0.022
r 24000_10000_M2 24000_12000_M2 0.022
r 24000_12000_M2 24000_14000_M2 0.022
r 24000_14000_M2 24000_16000_M2 0.022
r 24000_16000_M2 24000_18000_M2 0.022
r 24000_18000_M2 24000_20000_M2 0.022
r 24000_20000_M2 24000_22000_M2 0.022
r 24000_22000_M2 24000_24000_M2 0.022
r 24000_24000_M2 24000_26000_M2 0.022
r 24000_26000_M2 24000_28000_M2 0.022
r 24000_28000_M2 24000_30000_M2 0.022
r 24000_30000_M2 24000_32000_M2 0.022
r 24000_32000_M2 24000_34000_M2 0.022
r 24000_34000_M2 24000_36000_M2 0.022
r 24000_36000_M2 24000_38000_M2 0.022
r 24000_38000_M2 24000_40000_M2 0.022
r 24000_40000_M2 24000_42000_M2 0.022
r 24000_42000_M2 24000_44000_M2 0.022
r 24000_44000_M2 24000_46000_M2 0.022
r 24000_46000_M2 24000_48000_M2 0.022
r 24000_48000_M2 24000_50000_M2 0.022
r 24000_50000_M2 24000_52000_M2 0.022
r 24000_52000_M2 24000_54000_M2 0.022
r 24000_54000_M2 24000_56000_M2 0.022
r 24000_56000_M2 24000_58000_M2 0.022
r 24000_58000_M2 24000_60000_M2 0.022
r 24000_60000_M2 24000_62000_M2 0.022
r 24000_62000_M2 24000_64000_M2 0.022
r 24000_64000_M2 24000_66000_M2 0.022
r 24000_66000_M2 24000_68000_M2 0.022
r 24000_68000_M2 24000_70000_M2 0.022
r 24000_70000_M2 24000_72000_M2 0.022
r 24000_72000_M2 24000_74000_M2 0.022
r 24000_74000_M2 24000_76000_M2 0.022
r 24000_76000_M2 24000_78000_M2 0.022
r 24000_78000_M2 24000_80000_M2 0.022
r 24000_80000_M2 24000_82000_M2 0.022
r 24000_82000_M2 24000_84000_M2 0.022
r 24000_84000_M2 24000_86000_M2 0.022
r 24000_86000_M2 24000_88000_M2 0.022
r 24000_88000_M2 24000_90000_M2 0.022
r 24000_90000_M2 24000_92000_M2 0.022
r 24000_92000_M2 24000_94000_M2 0.022
r 24000_94000_M2 24000_96000_M2 0.022
r 24000_96000_M2 24000_98000_M2 0.022
r 24000_98000_M2 24000_100000_M2 0.022
r 26000_2000_M2 26000_4000_M2 0.022
r 26000_4000_M2 26000_6000_M2 0.022
r 26000_6000_M2 26000_8000_M2 0.022
r 26000_8000_M2 26000_10000_M2 0.022
r 26000_10000_M2 26000_12000_M2 0.022
r 26000_12000_M2 26000_14000_M2 0.022
r 26000_14000_M2 26000_16000_M2 0.022
r 26000_16000_M2 26000_18000_M2 0.022
r 26000_18000_M2 26000_20000_M2 0.022
r 26000_20000_M2 26000_22000_M2 0.022
r 26000_22000_M2 26000_24000_M2 0.022
r 26000_24000_M2 26000_26000_M2 0.022
r 26000_26000_M2 26000_28000_M2 0.022
r 26000_28000_M2 26000_30000_M2 0.022
r 26000_30000_M2 26000_32000_M2 0.022
r 26000_32000_M2 26000_34000_M2 0.022
r 26000_34000_M2 26000_36000_M2 0.022
r 26000_36000_M2 26000_38000_M2 0.022
r 26000_38000_M2 26000_40000_M2 0.022
r 26000_40000_M2 26000_42000_M2 0.022
r 26000_42000_M2 26000_44000_M2 0.022
r 26000_44000_M2 26000_46000_M2 0.022
r 26000_46000_M2 26000_48000_M2 0.022
r 26000_48000_M2 26000_50000_M2 0.022
r 26000_50000_M2 26000_52000_M2 0.022
r 26000_52000_M2 26000_54000_M2 0.022
r 26000_54000_M2 26000_56000_M2 0.022
r 26000_56000_M2 26000_58000_M2 0.022
r 26000_58000_M2 26000_60000_M2 0.022
r 26000_60000_M2 26000_62000_M2 0.022
r 26000_62000_M2 26000_64000_M2 0.022
r 26000_64000_M2 26000_66000_M2 0.022
r 26000_66000_M2 26000_68000_M2 0.022
r 26000_68000_M2 26000_70000_M2 0.022
r 26000_70000_M2 26000_72000_M2 0.022
r 26000_72000_M2 26000_74000_M2 0.022
r 26000_74000_M2 26000_76000_M2 0.022
r 26000_76000_M2 26000_78000_M2 0.022
r 26000_78000_M2 26000_80000_M2 0.022
r 26000_80000_M2 26000_82000_M2 0.022
r 26000_82000_M2 26000_84000_M2 0.022
r 26000_84000_M2 26000_86000_M2 0.022
r 26000_86000_M2 26000_88000_M2 0.022
r 26000_88000_M2 26000_90000_M2 0.022
r 26000_90000_M2 26000_92000_M2 0.022
r 26000_92000_M2 26000_94000_M2 0.022
r 26000_94000_M2 26000_96000_M2 0.022
r 26000_96000_M2 26000_98000_M2 0.022
r 26000_98000_M2 26000_100000_M2 0.022
r 28000_2000_M2 28000_4000_M2 0.022
r 28000_4000_M2 28000_6000_M2 0.022
r 28000_6000_M2 28000_8000_M2 0.022
r 28000_8000_M2 28000_10000_M2 0.022
r 28000_10000_M2 28000_12000_M2 0.022
r 28000_12000_M2 28000_14000_M2 0.022
r 28000_14000_M2 28000_16000_M2 0.022
r 28000_16000_M2 28000_18000_M2 0.022
r 28000_18000_M2 28000_20000_M2 0.022
r 28000_20000_M2 28000_22000_M2 0.022
r 28000_22000_M2 28000_24000_M2 0.022
r 28000_24000_M2 28000_26000_M2 0.022
r 28000_26000_M2 28000_28000_M2 0.022
r 28000_28000_M2 28000_30000_M2 0.022
r 28000_30000_M2 28000_32000_M2 0.022
r 28000_32000_M2 28000_34000_M2 0.022
r 28000_34000_M2 28000_36000_M2 0.022
r 28000_36000_M2 28000_38000_M2 0.022
r 28000_38000_M2 28000_40000_M2 0.022
r 28000_40000_M2 28000_42000_M2 0.022
r 28000_42000_M2 28000_44000_M2 0.022
r 28000_44000_M2 28000_46000_M2 0.022
r 28000_46000_M2 28000_48000_M2 0.022
r 28000_48000_M2 28000_50000_M2 0.022
r 28000_50000_M2 28000_52000_M2 0.022
r 28000_52000_M2 28000_54000_M2 0.022
r 28000_54000_M2 28000_56000_M2 0.022
r 28000_56000_M2 28000_58000_M2 0.022
r 28000_58000_M2 28000_60000_M2 0.022
r 28000_60000_M2 28000_62000_M2 0.022
r 28000_62000_M2 28000_64000_M2 0.022
r 28000_64000_M2 28000_66000_M2 0.022
r 28000_66000_M2 28000_68000_M2 0.022
r 28000_68000_M2 28000_70000_M2 0.022
r 28000_70000_M2 28000_72000_M2 0.022
r 28000_72000_M2 28000_74000_M2 0.022
r 28000_74000_M2 28000_76000_M2 0.022
r 28000_76000_M2 28000_78000_M2 0.022
r 28000_78000_M2 28000_80000_M2 0.022
r 28000_80000_M2 28000_82000_M2 0.022
r 28000_82000_M2 28000_84000_M2 0.022
r 28000_84000_M2 28000_86000_M2 0.022
r 28000_86000_M2 28000_88000_M2 0.022
r 28000_88000_M2 28000_90000_M2 0.022
r 28000_90000_M2 28000_92000_M2 0.022
r 28000_92000_M2 28000_94000_M2 0.022
r 28000_94000_M2 28000_96000_M2 0.022
r 28000_96000_M2 28000_98000_M2 0.022
r 28000_98000_M2 28000_100000_M2 0.022
r 30000_2000_M2 30000_4000_M2 0.022
r 30000_4000_M2 30000_6000_M2 0.022
r 30000_6000_M2 30000_8000_M2 0.022
r 30000_8000_M2 30000_10000_M2 0.022
r 30000_10000_M2 30000_12000_M2 0.022
r 30000_12000_M2 30000_14000_M2 0.022
r 30000_14000_M2 30000_16000_M2 0.022
r 30000_16000_M2 30000_18000_M2 0.022
r 30000_18000_M2 30000_20000_M2 0.022
r 30000_20000_M2 30000_22000_M2 0.022
r 30000_22000_M2 30000_24000_M2 0.022
r 30000_24000_M2 30000_26000_M2 0.022
r 30000_26000_M2 30000_28000_M2 0.022
r 30000_28000_M2 30000_30000_M2 0.022
r 30000_30000_M2 30000_32000_M2 0.022
r 30000_32000_M2 30000_34000_M2 0.022
r 30000_34000_M2 30000_36000_M2 0.022
r 30000_36000_M2 30000_38000_M2 0.022
r 30000_38000_M2 30000_40000_M2 0.022
r 30000_40000_M2 30000_42000_M2 0.022
r 30000_42000_M2 30000_44000_M2 0.022
r 30000_44000_M2 30000_46000_M2 0.022
r 30000_46000_M2 30000_48000_M2 0.022
r 30000_48000_M2 30000_50000_M2 0.022
r 30000_50000_M2 30000_52000_M2 0.022
r 30000_52000_M2 30000_54000_M2 0.022
r 30000_54000_M2 30000_56000_M2 0.022
r 30000_56000_M2 30000_58000_M2 0.022
r 30000_58000_M2 30000_60000_M2 0.022
r 30000_60000_M2 30000_62000_M2 0.022
r 30000_62000_M2 30000_64000_M2 0.022
r 30000_64000_M2 30000_66000_M2 0.022
r 30000_66000_M2 30000_68000_M2 0.022
r 30000_68000_M2 30000_70000_M2 0.022
r 30000_70000_M2 30000_72000_M2 0.022
r 30000_72000_M2 30000_74000_M2 0.022
r 30000_74000_M2 30000_76000_M2 0.022
r 30000_76000_M2 30000_78000_M2 0.022
r 30000_78000_M2 30000_80000_M2 0.022
r 30000_80000_M2 30000_82000_M2 0.022
r 30000_82000_M2 30000_84000_M2 0.022
r 30000_84000_M2 30000_86000_M2 0.022
r 30000_86000_M2 30000_88000_M2 0.022
r 30000_88000_M2 30000_90000_M2 0.022
r 30000_90000_M2 30000_92000_M2 0.022
r 30000_92000_M2 30000_94000_M2 0.022
r 30000_94000_M2 30000_96000_M2 0.022
r 30000_96000_M2 30000_98000_M2 0.022
r 30000_98000_M2 30000_100000_M2 0.022
r 32000_2000_M2 32000_4000_M2 0.022
r 32000_4000_M2 32000_6000_M2 0.022
r 32000_6000_M2 32000_8000_M2 0.022
r 32000_8000_M2 32000_10000_M2 0.022
r 32000_10000_M2 32000_12000_M2 0.022
r 32000_12000_M2 32000_14000_M2 0.022
r 32000_14000_M2 32000_16000_M2 0.022
r 32000_16000_M2 32000_18000_M2 0.022
r 32000_18000_M2 32000_20000_M2 0.022
r 32000_20000_M2 32000_22000_M2 0.022
r 32000_22000_M2 32000_24000_M2 0.022
r 32000_24000_M2 32000_26000_M2 0.022
r 32000_26000_M2 32000_28000_M2 0.022
r 32000_28000_M2 32000_30000_M2 0.022
r 32000_30000_M2 32000_32000_M2 0.022
r 32000_32000_M2 32000_34000_M2 0.022
r 32000_34000_M2 32000_36000_M2 0.022
r 32000_36000_M2 32000_38000_M2 0.022
r 32000_38000_M2 32000_40000_M2 0.022
r 32000_40000_M2 32000_42000_M2 0.022
r 32000_42000_M2 32000_44000_M2 0.022
r 32000_44000_M2 32000_46000_M2 0.022
r 32000_46000_M2 32000_48000_M2 0.022
r 32000_48000_M2 32000_50000_M2 0.022
r 32000_50000_M2 32000_52000_M2 0.022
r 32000_52000_M2 32000_54000_M2 0.022
r 32000_54000_M2 32000_56000_M2 0.022
r 32000_56000_M2 32000_58000_M2 0.022
r 32000_58000_M2 32000_60000_M2 0.022
r 32000_60000_M2 32000_62000_M2 0.022
r 32000_62000_M2 32000_64000_M2 0.022
r 32000_64000_M2 32000_66000_M2 0.022
r 32000_66000_M2 32000_68000_M2 0.022
r 32000_68000_M2 32000_70000_M2 0.022
r 32000_70000_M2 32000_72000_M2 0.022
r 32000_72000_M2 32000_74000_M2 0.022
r 32000_74000_M2 32000_76000_M2 0.022
r 32000_76000_M2 32000_78000_M2 0.022
r 32000_78000_M2 32000_80000_M2 0.022
r 32000_80000_M2 32000_82000_M2 0.022
r 32000_82000_M2 32000_84000_M2 0.022
r 32000_84000_M2 32000_86000_M2 0.022
r 32000_86000_M2 32000_88000_M2 0.022
r 32000_88000_M2 32000_90000_M2 0.022
r 32000_90000_M2 32000_92000_M2 0.022
r 32000_92000_M2 32000_94000_M2 0.022
r 32000_94000_M2 32000_96000_M2 0.022
r 32000_96000_M2 32000_98000_M2 0.022
r 32000_98000_M2 32000_100000_M2 0.022
r 34000_2000_M2 34000_4000_M2 0.022
r 34000_4000_M2 34000_6000_M2 0.022
r 34000_6000_M2 34000_8000_M2 0.022
r 34000_8000_M2 34000_10000_M2 0.022
r 34000_10000_M2 34000_12000_M2 0.022
r 34000_12000_M2 34000_14000_M2 0.022
r 34000_14000_M2 34000_16000_M2 0.022
r 34000_16000_M2 34000_18000_M2 0.022
r 34000_18000_M2 34000_20000_M2 0.022
r 34000_20000_M2 34000_22000_M2 0.022
r 34000_22000_M2 34000_24000_M2 0.022
r 34000_24000_M2 34000_26000_M2 0.022
r 34000_26000_M2 34000_28000_M2 0.022
r 34000_28000_M2 34000_30000_M2 0.022
r 34000_30000_M2 34000_32000_M2 0.022
r 34000_32000_M2 34000_34000_M2 0.022
r 34000_34000_M2 34000_36000_M2 0.022
r 34000_36000_M2 34000_38000_M2 0.022
r 34000_38000_M2 34000_40000_M2 0.022
r 34000_40000_M2 34000_42000_M2 0.022
r 34000_42000_M2 34000_44000_M2 0.022
r 34000_44000_M2 34000_46000_M2 0.022
r 34000_46000_M2 34000_48000_M2 0.022
r 34000_48000_M2 34000_50000_M2 0.022
r 34000_50000_M2 34000_52000_M2 0.022
r 34000_52000_M2 34000_54000_M2 0.022
r 34000_54000_M2 34000_56000_M2 0.022
r 34000_56000_M2 34000_58000_M2 0.022
r 34000_58000_M2 34000_60000_M2 0.022
r 34000_60000_M2 34000_62000_M2 0.022
r 34000_62000_M2 34000_64000_M2 0.022
r 34000_64000_M2 34000_66000_M2 0.022
r 34000_66000_M2 34000_68000_M2 0.022
r 34000_68000_M2 34000_70000_M2 0.022
r 34000_70000_M2 34000_72000_M2 0.022
r 34000_72000_M2 34000_74000_M2 0.022
r 34000_74000_M2 34000_76000_M2 0.022
r 34000_76000_M2 34000_78000_M2 0.022
r 34000_78000_M2 34000_80000_M2 0.022
r 34000_80000_M2 34000_82000_M2 0.022
r 34000_82000_M2 34000_84000_M2 0.022
r 34000_84000_M2 34000_86000_M2 0.022
r 34000_86000_M2 34000_88000_M2 0.022
r 34000_88000_M2 34000_90000_M2 0.022
r 34000_90000_M2 34000_92000_M2 0.022
r 34000_92000_M2 34000_94000_M2 0.022
r 34000_94000_M2 34000_96000_M2 0.022
r 34000_96000_M2 34000_98000_M2 0.022
r 34000_98000_M2 34000_100000_M2 0.022
r 36000_2000_M2 36000_4000_M2 0.022
r 36000_4000_M2 36000_6000_M2 0.022
r 36000_6000_M2 36000_8000_M2 0.022
r 36000_8000_M2 36000_10000_M2 0.022
r 36000_10000_M2 36000_12000_M2 0.022
r 36000_12000_M2 36000_14000_M2 0.022
r 36000_14000_M2 36000_16000_M2 0.022
r 36000_16000_M2 36000_18000_M2 0.022
r 36000_18000_M2 36000_20000_M2 0.022
r 36000_20000_M2 36000_22000_M2 0.022
r 36000_22000_M2 36000_24000_M2 0.022
r 36000_24000_M2 36000_26000_M2 0.022
r 36000_26000_M2 36000_28000_M2 0.022
r 36000_28000_M2 36000_30000_M2 0.022
r 36000_30000_M2 36000_32000_M2 0.022
r 36000_32000_M2 36000_34000_M2 0.022
r 36000_34000_M2 36000_36000_M2 0.022
r 36000_36000_M2 36000_38000_M2 0.022
r 36000_38000_M2 36000_40000_M2 0.022
r 36000_40000_M2 36000_42000_M2 0.022
r 36000_42000_M2 36000_44000_M2 0.022
r 36000_44000_M2 36000_46000_M2 0.022
r 36000_46000_M2 36000_48000_M2 0.022
r 36000_48000_M2 36000_50000_M2 0.022
r 36000_50000_M2 36000_52000_M2 0.022
r 36000_52000_M2 36000_54000_M2 0.022
r 36000_54000_M2 36000_56000_M2 0.022
r 36000_56000_M2 36000_58000_M2 0.022
r 36000_58000_M2 36000_60000_M2 0.022
r 36000_60000_M2 36000_62000_M2 0.022
r 36000_62000_M2 36000_64000_M2 0.022
r 36000_64000_M2 36000_66000_M2 0.022
r 36000_66000_M2 36000_68000_M2 0.022
r 36000_68000_M2 36000_70000_M2 0.022
r 36000_70000_M2 36000_72000_M2 0.022
r 36000_72000_M2 36000_74000_M2 0.022
r 36000_74000_M2 36000_76000_M2 0.022
r 36000_76000_M2 36000_78000_M2 0.022
r 36000_78000_M2 36000_80000_M2 0.022
r 36000_80000_M2 36000_82000_M2 0.022
r 36000_82000_M2 36000_84000_M2 0.022
r 36000_84000_M2 36000_86000_M2 0.022
r 36000_86000_M2 36000_88000_M2 0.022
r 36000_88000_M2 36000_90000_M2 0.022
r 36000_90000_M2 36000_92000_M2 0.022
r 36000_92000_M2 36000_94000_M2 0.022
r 36000_94000_M2 36000_96000_M2 0.022
r 36000_96000_M2 36000_98000_M2 0.022
r 36000_98000_M2 36000_100000_M2 0.022
r 38000_2000_M2 38000_4000_M2 0.022
r 38000_4000_M2 38000_6000_M2 0.022
r 38000_6000_M2 38000_8000_M2 0.022
r 38000_8000_M2 38000_10000_M2 0.022
r 38000_10000_M2 38000_12000_M2 0.022
r 38000_12000_M2 38000_14000_M2 0.022
r 38000_14000_M2 38000_16000_M2 0.022
r 38000_16000_M2 38000_18000_M2 0.022
r 38000_18000_M2 38000_20000_M2 0.022
r 38000_20000_M2 38000_22000_M2 0.022
r 38000_22000_M2 38000_24000_M2 0.022
r 38000_24000_M2 38000_26000_M2 0.022
r 38000_26000_M2 38000_28000_M2 0.022
r 38000_28000_M2 38000_30000_M2 0.022
r 38000_30000_M2 38000_32000_M2 0.022
r 38000_32000_M2 38000_34000_M2 0.022
r 38000_34000_M2 38000_36000_M2 0.022
r 38000_36000_M2 38000_38000_M2 0.022
r 38000_38000_M2 38000_40000_M2 0.022
r 38000_40000_M2 38000_42000_M2 0.022
r 38000_42000_M2 38000_44000_M2 0.022
r 38000_44000_M2 38000_46000_M2 0.022
r 38000_46000_M2 38000_48000_M2 0.022
r 38000_48000_M2 38000_50000_M2 0.022
r 38000_50000_M2 38000_52000_M2 0.022
r 38000_52000_M2 38000_54000_M2 0.022
r 38000_54000_M2 38000_56000_M2 0.022
r 38000_56000_M2 38000_58000_M2 0.022
r 38000_58000_M2 38000_60000_M2 0.022
r 38000_60000_M2 38000_62000_M2 0.022
r 38000_62000_M2 38000_64000_M2 0.022
r 38000_64000_M2 38000_66000_M2 0.022
r 38000_66000_M2 38000_68000_M2 0.022
r 38000_68000_M2 38000_70000_M2 0.022
r 38000_70000_M2 38000_72000_M2 0.022
r 38000_72000_M2 38000_74000_M2 0.022
r 38000_74000_M2 38000_76000_M2 0.022
r 38000_76000_M2 38000_78000_M2 0.022
r 38000_78000_M2 38000_80000_M2 0.022
r 38000_80000_M2 38000_82000_M2 0.022
r 38000_82000_M2 38000_84000_M2 0.022
r 38000_84000_M2 38000_86000_M2 0.022
r 38000_86000_M2 38000_88000_M2 0.022
r 38000_88000_M2 38000_90000_M2 0.022
r 38000_90000_M2 38000_92000_M2 0.022
r 38000_92000_M2 38000_94000_M2 0.022
r 38000_94000_M2 38000_96000_M2 0.022
r 38000_96000_M2 38000_98000_M2 0.022
r 38000_98000_M2 38000_100000_M2 0.022
r 40000_2000_M2 40000_4000_M2 0.022
r 40000_4000_M2 40000_6000_M2 0.022
r 40000_6000_M2 40000_8000_M2 0.022
r 40000_8000_M2 40000_10000_M2 0.022
r 40000_10000_M2 40000_12000_M2 0.022
r 40000_12000_M2 40000_14000_M2 0.022
r 40000_14000_M2 40000_16000_M2 0.022
r 40000_16000_M2 40000_18000_M2 0.022
r 40000_18000_M2 40000_20000_M2 0.022
r 40000_20000_M2 40000_22000_M2 0.022
r 40000_22000_M2 40000_24000_M2 0.022
r 40000_24000_M2 40000_26000_M2 0.022
r 40000_26000_M2 40000_28000_M2 0.022
r 40000_28000_M2 40000_30000_M2 0.022
r 40000_30000_M2 40000_32000_M2 0.022
r 40000_32000_M2 40000_34000_M2 0.022
r 40000_34000_M2 40000_36000_M2 0.022
r 40000_36000_M2 40000_38000_M2 0.022
r 40000_38000_M2 40000_40000_M2 0.022
r 40000_40000_M2 40000_42000_M2 0.022
r 40000_42000_M2 40000_44000_M2 0.022
r 40000_44000_M2 40000_46000_M2 0.022
r 40000_46000_M2 40000_48000_M2 0.022
r 40000_48000_M2 40000_50000_M2 0.022
r 40000_50000_M2 40000_52000_M2 0.022
r 40000_52000_M2 40000_54000_M2 0.022
r 40000_54000_M2 40000_56000_M2 0.022
r 40000_56000_M2 40000_58000_M2 0.022
r 40000_58000_M2 40000_60000_M2 0.022
r 40000_60000_M2 40000_62000_M2 0.022
r 40000_62000_M2 40000_64000_M2 0.022
r 40000_64000_M2 40000_66000_M2 0.022
r 40000_66000_M2 40000_68000_M2 0.022
r 40000_68000_M2 40000_70000_M2 0.022
r 40000_70000_M2 40000_72000_M2 0.022
r 40000_72000_M2 40000_74000_M2 0.022
r 40000_74000_M2 40000_76000_M2 0.022
r 40000_76000_M2 40000_78000_M2 0.022
r 40000_78000_M2 40000_80000_M2 0.022
r 40000_80000_M2 40000_82000_M2 0.022
r 40000_82000_M2 40000_84000_M2 0.022
r 40000_84000_M2 40000_86000_M2 0.022
r 40000_86000_M2 40000_88000_M2 0.022
r 40000_88000_M2 40000_90000_M2 0.022
r 40000_90000_M2 40000_92000_M2 0.022
r 40000_92000_M2 40000_94000_M2 0.022
r 40000_94000_M2 40000_96000_M2 0.022
r 40000_96000_M2 40000_98000_M2 0.022
r 40000_98000_M2 40000_100000_M2 0.022
r 42000_2000_M2 42000_4000_M2 0.022
r 42000_4000_M2 42000_6000_M2 0.022
r 42000_6000_M2 42000_8000_M2 0.022
r 42000_8000_M2 42000_10000_M2 0.022
r 42000_10000_M2 42000_12000_M2 0.022
r 42000_12000_M2 42000_14000_M2 0.022
r 42000_14000_M2 42000_16000_M2 0.022
r 42000_16000_M2 42000_18000_M2 0.022
r 42000_18000_M2 42000_20000_M2 0.022
r 42000_20000_M2 42000_22000_M2 0.022
r 42000_22000_M2 42000_24000_M2 0.022
r 42000_24000_M2 42000_26000_M2 0.022
r 42000_26000_M2 42000_28000_M2 0.022
r 42000_28000_M2 42000_30000_M2 0.022
r 42000_30000_M2 42000_32000_M2 0.022
r 42000_32000_M2 42000_34000_M2 0.022
r 42000_34000_M2 42000_36000_M2 0.022
r 42000_36000_M2 42000_38000_M2 0.022
r 42000_38000_M2 42000_40000_M2 0.022
r 42000_40000_M2 42000_42000_M2 0.022
r 42000_42000_M2 42000_44000_M2 0.022
r 42000_44000_M2 42000_46000_M2 0.022
r 42000_46000_M2 42000_48000_M2 0.022
r 42000_48000_M2 42000_50000_M2 0.022
r 42000_50000_M2 42000_52000_M2 0.022
r 42000_52000_M2 42000_54000_M2 0.022
r 42000_54000_M2 42000_56000_M2 0.022
r 42000_56000_M2 42000_58000_M2 0.022
r 42000_58000_M2 42000_60000_M2 0.022
r 42000_60000_M2 42000_62000_M2 0.022
r 42000_62000_M2 42000_64000_M2 0.022
r 42000_64000_M2 42000_66000_M2 0.022
r 42000_66000_M2 42000_68000_M2 0.022
r 42000_68000_M2 42000_70000_M2 0.022
r 42000_70000_M2 42000_72000_M2 0.022
r 42000_72000_M2 42000_74000_M2 0.022
r 42000_74000_M2 42000_76000_M2 0.022
r 42000_76000_M2 42000_78000_M2 0.022
r 42000_78000_M2 42000_80000_M2 0.022
r 42000_80000_M2 42000_82000_M2 0.022
r 42000_82000_M2 42000_84000_M2 0.022
r 42000_84000_M2 42000_86000_M2 0.022
r 42000_86000_M2 42000_88000_M2 0.022
r 42000_88000_M2 42000_90000_M2 0.022
r 42000_90000_M2 42000_92000_M2 0.022
r 42000_92000_M2 42000_94000_M2 0.022
r 42000_94000_M2 42000_96000_M2 0.022
r 42000_96000_M2 42000_98000_M2 0.022
r 42000_98000_M2 42000_100000_M2 0.022
r 44000_2000_M2 44000_4000_M2 0.022
r 44000_4000_M2 44000_6000_M2 0.022
r 44000_6000_M2 44000_8000_M2 0.022
r 44000_8000_M2 44000_10000_M2 0.022
r 44000_10000_M2 44000_12000_M2 0.022
r 44000_12000_M2 44000_14000_M2 0.022
r 44000_14000_M2 44000_16000_M2 0.022
r 44000_16000_M2 44000_18000_M2 0.022
r 44000_18000_M2 44000_20000_M2 0.022
r 44000_20000_M2 44000_22000_M2 0.022
r 44000_22000_M2 44000_24000_M2 0.022
r 44000_24000_M2 44000_26000_M2 0.022
r 44000_26000_M2 44000_28000_M2 0.022
r 44000_28000_M2 44000_30000_M2 0.022
r 44000_30000_M2 44000_32000_M2 0.022
r 44000_32000_M2 44000_34000_M2 0.022
r 44000_34000_M2 44000_36000_M2 0.022
r 44000_36000_M2 44000_38000_M2 0.022
r 44000_38000_M2 44000_40000_M2 0.022
r 44000_40000_M2 44000_42000_M2 0.022
r 44000_42000_M2 44000_44000_M2 0.022
r 44000_44000_M2 44000_46000_M2 0.022
r 44000_46000_M2 44000_48000_M2 0.022
r 44000_48000_M2 44000_50000_M2 0.022
r 44000_50000_M2 44000_52000_M2 0.022
r 44000_52000_M2 44000_54000_M2 0.022
r 44000_54000_M2 44000_56000_M2 0.022
r 44000_56000_M2 44000_58000_M2 0.022
r 44000_58000_M2 44000_60000_M2 0.022
r 44000_60000_M2 44000_62000_M2 0.022
r 44000_62000_M2 44000_64000_M2 0.022
r 44000_64000_M2 44000_66000_M2 0.022
r 44000_66000_M2 44000_68000_M2 0.022
r 44000_68000_M2 44000_70000_M2 0.022
r 44000_70000_M2 44000_72000_M2 0.022
r 44000_72000_M2 44000_74000_M2 0.022
r 44000_74000_M2 44000_76000_M2 0.022
r 44000_76000_M2 44000_78000_M2 0.022
r 44000_78000_M2 44000_80000_M2 0.022
r 44000_80000_M2 44000_82000_M2 0.022
r 44000_82000_M2 44000_84000_M2 0.022
r 44000_84000_M2 44000_86000_M2 0.022
r 44000_86000_M2 44000_88000_M2 0.022
r 44000_88000_M2 44000_90000_M2 0.022
r 44000_90000_M2 44000_92000_M2 0.022
r 44000_92000_M2 44000_94000_M2 0.022
r 44000_94000_M2 44000_96000_M2 0.022
r 44000_96000_M2 44000_98000_M2 0.022
r 44000_98000_M2 44000_100000_M2 0.022
r 46000_2000_M2 46000_4000_M2 0.022
r 46000_4000_M2 46000_6000_M2 0.022
r 46000_6000_M2 46000_8000_M2 0.022
r 46000_8000_M2 46000_10000_M2 0.022
r 46000_10000_M2 46000_12000_M2 0.022
r 46000_12000_M2 46000_14000_M2 0.022
r 46000_14000_M2 46000_16000_M2 0.022
r 46000_16000_M2 46000_18000_M2 0.022
r 46000_18000_M2 46000_20000_M2 0.022
r 46000_20000_M2 46000_22000_M2 0.022
r 46000_22000_M2 46000_24000_M2 0.022
r 46000_24000_M2 46000_26000_M2 0.022
r 46000_26000_M2 46000_28000_M2 0.022
r 46000_28000_M2 46000_30000_M2 0.022
r 46000_30000_M2 46000_32000_M2 0.022
r 46000_32000_M2 46000_34000_M2 0.022
r 46000_34000_M2 46000_36000_M2 0.022
r 46000_36000_M2 46000_38000_M2 0.022
r 46000_38000_M2 46000_40000_M2 0.022
r 46000_40000_M2 46000_42000_M2 0.022
r 46000_42000_M2 46000_44000_M2 0.022
r 46000_44000_M2 46000_46000_M2 0.022
r 46000_46000_M2 46000_48000_M2 0.022
r 46000_48000_M2 46000_50000_M2 0.022
r 46000_50000_M2 46000_52000_M2 0.022
r 46000_52000_M2 46000_54000_M2 0.022
r 46000_54000_M2 46000_56000_M2 0.022
r 46000_56000_M2 46000_58000_M2 0.022
r 46000_58000_M2 46000_60000_M2 0.022
r 46000_60000_M2 46000_62000_M2 0.022
r 46000_62000_M2 46000_64000_M2 0.022
r 46000_64000_M2 46000_66000_M2 0.022
r 46000_66000_M2 46000_68000_M2 0.022
r 46000_68000_M2 46000_70000_M2 0.022
r 46000_70000_M2 46000_72000_M2 0.022
r 46000_72000_M2 46000_74000_M2 0.022
r 46000_74000_M2 46000_76000_M2 0.022
r 46000_76000_M2 46000_78000_M2 0.022
r 46000_78000_M2 46000_80000_M2 0.022
r 46000_80000_M2 46000_82000_M2 0.022
r 46000_82000_M2 46000_84000_M2 0.022
r 46000_84000_M2 46000_86000_M2 0.022
r 46000_86000_M2 46000_88000_M2 0.022
r 46000_88000_M2 46000_90000_M2 0.022
r 46000_90000_M2 46000_92000_M2 0.022
r 46000_92000_M2 46000_94000_M2 0.022
r 46000_94000_M2 46000_96000_M2 0.022
r 46000_96000_M2 46000_98000_M2 0.022
r 46000_98000_M2 46000_100000_M2 0.022
r 48000_2000_M2 48000_4000_M2 0.022
r 48000_4000_M2 48000_6000_M2 0.022
r 48000_6000_M2 48000_8000_M2 0.022
r 48000_8000_M2 48000_10000_M2 0.022
r 48000_10000_M2 48000_12000_M2 0.022
r 48000_12000_M2 48000_14000_M2 0.022
r 48000_14000_M2 48000_16000_M2 0.022
r 48000_16000_M2 48000_18000_M2 0.022
r 48000_18000_M2 48000_20000_M2 0.022
r 48000_20000_M2 48000_22000_M2 0.022
r 48000_22000_M2 48000_24000_M2 0.022
r 48000_24000_M2 48000_26000_M2 0.022
r 48000_26000_M2 48000_28000_M2 0.022
r 48000_28000_M2 48000_30000_M2 0.022
r 48000_30000_M2 48000_32000_M2 0.022
r 48000_32000_M2 48000_34000_M2 0.022
r 48000_34000_M2 48000_36000_M2 0.022
r 48000_36000_M2 48000_38000_M2 0.022
r 48000_38000_M2 48000_40000_M2 0.022
r 48000_40000_M2 48000_42000_M2 0.022
r 48000_42000_M2 48000_44000_M2 0.022
r 48000_44000_M2 48000_46000_M2 0.022
r 48000_46000_M2 48000_48000_M2 0.022
r 48000_48000_M2 48000_50000_M2 0.022
r 48000_50000_M2 48000_52000_M2 0.022
r 48000_52000_M2 48000_54000_M2 0.022
r 48000_54000_M2 48000_56000_M2 0.022
r 48000_56000_M2 48000_58000_M2 0.022
r 48000_58000_M2 48000_60000_M2 0.022
r 48000_60000_M2 48000_62000_M2 0.022
r 48000_62000_M2 48000_64000_M2 0.022
r 48000_64000_M2 48000_66000_M2 0.022
r 48000_66000_M2 48000_68000_M2 0.022
r 48000_68000_M2 48000_70000_M2 0.022
r 48000_70000_M2 48000_72000_M2 0.022
r 48000_72000_M2 48000_74000_M2 0.022
r 48000_74000_M2 48000_76000_M2 0.022
r 48000_76000_M2 48000_78000_M2 0.022
r 48000_78000_M2 48000_80000_M2 0.022
r 48000_80000_M2 48000_82000_M2 0.022
r 48000_82000_M2 48000_84000_M2 0.022
r 48000_84000_M2 48000_86000_M2 0.022
r 48000_86000_M2 48000_88000_M2 0.022
r 48000_88000_M2 48000_90000_M2 0.022
r 48000_90000_M2 48000_92000_M2 0.022
r 48000_92000_M2 48000_94000_M2 0.022
r 48000_94000_M2 48000_96000_M2 0.022
r 48000_96000_M2 48000_98000_M2 0.022
r 48000_98000_M2 48000_100000_M2 0.022
r 50000_2000_M2 50000_4000_M2 0.022
r 50000_4000_M2 50000_6000_M2 0.022
r 50000_6000_M2 50000_8000_M2 0.022
r 50000_8000_M2 50000_10000_M2 0.022
r 50000_10000_M2 50000_12000_M2 0.022
r 50000_12000_M2 50000_14000_M2 0.022
r 50000_14000_M2 50000_16000_M2 0.022
r 50000_16000_M2 50000_18000_M2 0.022
r 50000_18000_M2 50000_20000_M2 0.022
r 50000_20000_M2 50000_22000_M2 0.022
r 50000_22000_M2 50000_24000_M2 0.022
r 50000_24000_M2 50000_26000_M2 0.022
r 50000_26000_M2 50000_28000_M2 0.022
r 50000_28000_M2 50000_30000_M2 0.022
r 50000_30000_M2 50000_32000_M2 0.022
r 50000_32000_M2 50000_34000_M2 0.022
r 50000_34000_M2 50000_36000_M2 0.022
r 50000_36000_M2 50000_38000_M2 0.022
r 50000_38000_M2 50000_40000_M2 0.022
r 50000_40000_M2 50000_42000_M2 0.022
r 50000_42000_M2 50000_44000_M2 0.022
r 50000_44000_M2 50000_46000_M2 0.022
r 50000_46000_M2 50000_48000_M2 0.022
r 50000_48000_M2 50000_50000_M2 0.022
r 50000_50000_M2 50000_52000_M2 0.022
r 50000_52000_M2 50000_54000_M2 0.022
r 50000_54000_M2 50000_56000_M2 0.022
r 50000_56000_M2 50000_58000_M2 0.022
r 50000_58000_M2 50000_60000_M2 0.022
r 50000_60000_M2 50000_62000_M2 0.022
r 50000_62000_M2 50000_64000_M2 0.022
r 50000_64000_M2 50000_66000_M2 0.022
r 50000_66000_M2 50000_68000_M2 0.022
r 50000_68000_M2 50000_70000_M2 0.022
r 50000_70000_M2 50000_72000_M2 0.022
r 50000_72000_M2 50000_74000_M2 0.022
r 50000_74000_M2 50000_76000_M2 0.022
r 50000_76000_M2 50000_78000_M2 0.022
r 50000_78000_M2 50000_80000_M2 0.022
r 50000_80000_M2 50000_82000_M2 0.022
r 50000_82000_M2 50000_84000_M2 0.022
r 50000_84000_M2 50000_86000_M2 0.022
r 50000_86000_M2 50000_88000_M2 0.022
r 50000_88000_M2 50000_90000_M2 0.022
r 50000_90000_M2 50000_92000_M2 0.022
r 50000_92000_M2 50000_94000_M2 0.022
r 50000_94000_M2 50000_96000_M2 0.022
r 50000_96000_M2 50000_98000_M2 0.022
r 50000_98000_M2 50000_100000_M2 0.022
r 52000_2000_M2 52000_4000_M2 0.022
r 52000_4000_M2 52000_6000_M2 0.022
r 52000_6000_M2 52000_8000_M2 0.022
r 52000_8000_M2 52000_10000_M2 0.022
r 52000_10000_M2 52000_12000_M2 0.022
r 52000_12000_M2 52000_14000_M2 0.022
r 52000_14000_M2 52000_16000_M2 0.022
r 52000_16000_M2 52000_18000_M2 0.022
r 52000_18000_M2 52000_20000_M2 0.022
r 52000_20000_M2 52000_22000_M2 0.022
r 52000_22000_M2 52000_24000_M2 0.022
r 52000_24000_M2 52000_26000_M2 0.022
r 52000_26000_M2 52000_28000_M2 0.022
r 52000_28000_M2 52000_30000_M2 0.022
r 52000_30000_M2 52000_32000_M2 0.022
r 52000_32000_M2 52000_34000_M2 0.022
r 52000_34000_M2 52000_36000_M2 0.022
r 52000_36000_M2 52000_38000_M2 0.022
r 52000_38000_M2 52000_40000_M2 0.022
r 52000_40000_M2 52000_42000_M2 0.022
r 52000_42000_M2 52000_44000_M2 0.022
r 52000_44000_M2 52000_46000_M2 0.022
r 52000_46000_M2 52000_48000_M2 0.022
r 52000_48000_M2 52000_50000_M2 0.022
r 52000_50000_M2 52000_52000_M2 0.022
r 52000_52000_M2 52000_54000_M2 0.022
r 52000_54000_M2 52000_56000_M2 0.022
r 52000_56000_M2 52000_58000_M2 0.022
r 52000_58000_M2 52000_60000_M2 0.022
r 52000_60000_M2 52000_62000_M2 0.022
r 52000_62000_M2 52000_64000_M2 0.022
r 52000_64000_M2 52000_66000_M2 0.022
r 52000_66000_M2 52000_68000_M2 0.022
r 52000_68000_M2 52000_70000_M2 0.022
r 52000_70000_M2 52000_72000_M2 0.022
r 52000_72000_M2 52000_74000_M2 0.022
r 52000_74000_M2 52000_76000_M2 0.022
r 52000_76000_M2 52000_78000_M2 0.022
r 52000_78000_M2 52000_80000_M2 0.022
r 52000_80000_M2 52000_82000_M2 0.022
r 52000_82000_M2 52000_84000_M2 0.022
r 52000_84000_M2 52000_86000_M2 0.022
r 52000_86000_M2 52000_88000_M2 0.022
r 52000_88000_M2 52000_90000_M2 0.022
r 52000_90000_M2 52000_92000_M2 0.022
r 52000_92000_M2 52000_94000_M2 0.022
r 52000_94000_M2 52000_96000_M2 0.022
r 52000_96000_M2 52000_98000_M2 0.022
r 52000_98000_M2 52000_100000_M2 0.022
r 54000_2000_M2 54000_4000_M2 0.022
r 54000_4000_M2 54000_6000_M2 0.022
r 54000_6000_M2 54000_8000_M2 0.022
r 54000_8000_M2 54000_10000_M2 0.022
r 54000_10000_M2 54000_12000_M2 0.022
r 54000_12000_M2 54000_14000_M2 0.022
r 54000_14000_M2 54000_16000_M2 0.022
r 54000_16000_M2 54000_18000_M2 0.022
r 54000_18000_M2 54000_20000_M2 0.022
r 54000_20000_M2 54000_22000_M2 0.022
r 54000_22000_M2 54000_24000_M2 0.022
r 54000_24000_M2 54000_26000_M2 0.022
r 54000_26000_M2 54000_28000_M2 0.022
r 54000_28000_M2 54000_30000_M2 0.022
r 54000_30000_M2 54000_32000_M2 0.022
r 54000_32000_M2 54000_34000_M2 0.022
r 54000_34000_M2 54000_36000_M2 0.022
r 54000_36000_M2 54000_38000_M2 0.022
r 54000_38000_M2 54000_40000_M2 0.022
r 54000_40000_M2 54000_42000_M2 0.022
r 54000_42000_M2 54000_44000_M2 0.022
r 54000_44000_M2 54000_46000_M2 0.022
r 54000_46000_M2 54000_48000_M2 0.022
r 54000_48000_M2 54000_50000_M2 0.022
r 54000_50000_M2 54000_52000_M2 0.022
r 54000_52000_M2 54000_54000_M2 0.022
r 54000_54000_M2 54000_56000_M2 0.022
r 54000_56000_M2 54000_58000_M2 0.022
r 54000_58000_M2 54000_60000_M2 0.022
r 54000_60000_M2 54000_62000_M2 0.022
r 54000_62000_M2 54000_64000_M2 0.022
r 54000_64000_M2 54000_66000_M2 0.022
r 54000_66000_M2 54000_68000_M2 0.022
r 54000_68000_M2 54000_70000_M2 0.022
r 54000_70000_M2 54000_72000_M2 0.022
r 54000_72000_M2 54000_74000_M2 0.022
r 54000_74000_M2 54000_76000_M2 0.022
r 54000_76000_M2 54000_78000_M2 0.022
r 54000_78000_M2 54000_80000_M2 0.022
r 54000_80000_M2 54000_82000_M2 0.022
r 54000_82000_M2 54000_84000_M2 0.022
r 54000_84000_M2 54000_86000_M2 0.022
r 54000_86000_M2 54000_88000_M2 0.022
r 54000_88000_M2 54000_90000_M2 0.022
r 54000_90000_M2 54000_92000_M2 0.022
r 54000_92000_M2 54000_94000_M2 0.022
r 54000_94000_M2 54000_96000_M2 0.022
r 54000_96000_M2 54000_98000_M2 0.022
r 54000_98000_M2 54000_100000_M2 0.022
r 56000_2000_M2 56000_4000_M2 0.022
r 56000_4000_M2 56000_6000_M2 0.022
r 56000_6000_M2 56000_8000_M2 0.022
r 56000_8000_M2 56000_10000_M2 0.022
r 56000_10000_M2 56000_12000_M2 0.022
r 56000_12000_M2 56000_14000_M2 0.022
r 56000_14000_M2 56000_16000_M2 0.022
r 56000_16000_M2 56000_18000_M2 0.022
r 56000_18000_M2 56000_20000_M2 0.022
r 56000_20000_M2 56000_22000_M2 0.022
r 56000_22000_M2 56000_24000_M2 0.022
r 56000_24000_M2 56000_26000_M2 0.022
r 56000_26000_M2 56000_28000_M2 0.022
r 56000_28000_M2 56000_30000_M2 0.022
r 56000_30000_M2 56000_32000_M2 0.022
r 56000_32000_M2 56000_34000_M2 0.022
r 56000_34000_M2 56000_36000_M2 0.022
r 56000_36000_M2 56000_38000_M2 0.022
r 56000_38000_M2 56000_40000_M2 0.022
r 56000_40000_M2 56000_42000_M2 0.022
r 56000_42000_M2 56000_44000_M2 0.022
r 56000_44000_M2 56000_46000_M2 0.022
r 56000_46000_M2 56000_48000_M2 0.022
r 56000_48000_M2 56000_50000_M2 0.022
r 56000_50000_M2 56000_52000_M2 0.022
r 56000_52000_M2 56000_54000_M2 0.022
r 56000_54000_M2 56000_56000_M2 0.022
r 56000_56000_M2 56000_58000_M2 0.022
r 56000_58000_M2 56000_60000_M2 0.022
r 56000_60000_M2 56000_62000_M2 0.022
r 56000_62000_M2 56000_64000_M2 0.022
r 56000_64000_M2 56000_66000_M2 0.022
r 56000_66000_M2 56000_68000_M2 0.022
r 56000_68000_M2 56000_70000_M2 0.022
r 56000_70000_M2 56000_72000_M2 0.022
r 56000_72000_M2 56000_74000_M2 0.022
r 56000_74000_M2 56000_76000_M2 0.022
r 56000_76000_M2 56000_78000_M2 0.022
r 56000_78000_M2 56000_80000_M2 0.022
r 56000_80000_M2 56000_82000_M2 0.022
r 56000_82000_M2 56000_84000_M2 0.022
r 56000_84000_M2 56000_86000_M2 0.022
r 56000_86000_M2 56000_88000_M2 0.022
r 56000_88000_M2 56000_90000_M2 0.022
r 56000_90000_M2 56000_92000_M2 0.022
r 56000_92000_M2 56000_94000_M2 0.022
r 56000_94000_M2 56000_96000_M2 0.022
r 56000_96000_M2 56000_98000_M2 0.022
r 56000_98000_M2 56000_100000_M2 0.022
r 58000_2000_M2 58000_4000_M2 0.022
r 58000_4000_M2 58000_6000_M2 0.022
r 58000_6000_M2 58000_8000_M2 0.022
r 58000_8000_M2 58000_10000_M2 0.022
r 58000_10000_M2 58000_12000_M2 0.022
r 58000_12000_M2 58000_14000_M2 0.022
r 58000_14000_M2 58000_16000_M2 0.022
r 58000_16000_M2 58000_18000_M2 0.022
r 58000_18000_M2 58000_20000_M2 0.022
r 58000_20000_M2 58000_22000_M2 0.022
r 58000_22000_M2 58000_24000_M2 0.022
r 58000_24000_M2 58000_26000_M2 0.022
r 58000_26000_M2 58000_28000_M2 0.022
r 58000_28000_M2 58000_30000_M2 0.022
r 58000_30000_M2 58000_32000_M2 0.022
r 58000_32000_M2 58000_34000_M2 0.022
r 58000_34000_M2 58000_36000_M2 0.022
r 58000_36000_M2 58000_38000_M2 0.022
r 58000_38000_M2 58000_40000_M2 0.022
r 58000_40000_M2 58000_42000_M2 0.022
r 58000_42000_M2 58000_44000_M2 0.022
r 58000_44000_M2 58000_46000_M2 0.022
r 58000_46000_M2 58000_48000_M2 0.022
r 58000_48000_M2 58000_50000_M2 0.022
r 58000_50000_M2 58000_52000_M2 0.022
r 58000_52000_M2 58000_54000_M2 0.022
r 58000_54000_M2 58000_56000_M2 0.022
r 58000_56000_M2 58000_58000_M2 0.022
r 58000_58000_M2 58000_60000_M2 0.022
r 58000_60000_M2 58000_62000_M2 0.022
r 58000_62000_M2 58000_64000_M2 0.022
r 58000_64000_M2 58000_66000_M2 0.022
r 58000_66000_M2 58000_68000_M2 0.022
r 58000_68000_M2 58000_70000_M2 0.022
r 58000_70000_M2 58000_72000_M2 0.022
r 58000_72000_M2 58000_74000_M2 0.022
r 58000_74000_M2 58000_76000_M2 0.022
r 58000_76000_M2 58000_78000_M2 0.022
r 58000_78000_M2 58000_80000_M2 0.022
r 58000_80000_M2 58000_82000_M2 0.022
r 58000_82000_M2 58000_84000_M2 0.022
r 58000_84000_M2 58000_86000_M2 0.022
r 58000_86000_M2 58000_88000_M2 0.022
r 58000_88000_M2 58000_90000_M2 0.022
r 58000_90000_M2 58000_92000_M2 0.022
r 58000_92000_M2 58000_94000_M2 0.022
r 58000_94000_M2 58000_96000_M2 0.022
r 58000_96000_M2 58000_98000_M2 0.022
r 58000_98000_M2 58000_100000_M2 0.022
r 60000_2000_M2 60000_4000_M2 0.022
r 60000_4000_M2 60000_6000_M2 0.022
r 60000_6000_M2 60000_8000_M2 0.022
r 60000_8000_M2 60000_10000_M2 0.022
r 60000_10000_M2 60000_12000_M2 0.022
r 60000_12000_M2 60000_14000_M2 0.022
r 60000_14000_M2 60000_16000_M2 0.022
r 60000_16000_M2 60000_18000_M2 0.022
r 60000_18000_M2 60000_20000_M2 0.022
r 60000_20000_M2 60000_22000_M2 0.022
r 60000_22000_M2 60000_24000_M2 0.022
r 60000_24000_M2 60000_26000_M2 0.022
r 60000_26000_M2 60000_28000_M2 0.022
r 60000_28000_M2 60000_30000_M2 0.022
r 60000_30000_M2 60000_32000_M2 0.022
r 60000_32000_M2 60000_34000_M2 0.022
r 60000_34000_M2 60000_36000_M2 0.022
r 60000_36000_M2 60000_38000_M2 0.022
r 60000_38000_M2 60000_40000_M2 0.022
r 60000_40000_M2 60000_42000_M2 0.022
r 60000_42000_M2 60000_44000_M2 0.022
r 60000_44000_M2 60000_46000_M2 0.022
r 60000_46000_M2 60000_48000_M2 0.022
r 60000_48000_M2 60000_50000_M2 0.022
r 60000_50000_M2 60000_52000_M2 0.022
r 60000_52000_M2 60000_54000_M2 0.022
r 60000_54000_M2 60000_56000_M2 0.022
r 60000_56000_M2 60000_58000_M2 0.022
r 60000_58000_M2 60000_60000_M2 0.022
r 60000_60000_M2 60000_62000_M2 0.022
r 60000_62000_M2 60000_64000_M2 0.022
r 60000_64000_M2 60000_66000_M2 0.022
r 60000_66000_M2 60000_68000_M2 0.022
r 60000_68000_M2 60000_70000_M2 0.022
r 60000_70000_M2 60000_72000_M2 0.022
r 60000_72000_M2 60000_74000_M2 0.022
r 60000_74000_M2 60000_76000_M2 0.022
r 60000_76000_M2 60000_78000_M2 0.022
r 60000_78000_M2 60000_80000_M2 0.022
r 60000_80000_M2 60000_82000_M2 0.022
r 60000_82000_M2 60000_84000_M2 0.022
r 60000_84000_M2 60000_86000_M2 0.022
r 60000_86000_M2 60000_88000_M2 0.022
r 60000_88000_M2 60000_90000_M2 0.022
r 60000_90000_M2 60000_92000_M2 0.022
r 60000_92000_M2 60000_94000_M2 0.022
r 60000_94000_M2 60000_96000_M2 0.022
r 60000_96000_M2 60000_98000_M2 0.022
r 60000_98000_M2 60000_100000_M2 0.022
r 62000_2000_M2 62000_4000_M2 0.022
r 62000_4000_M2 62000_6000_M2 0.022
r 62000_6000_M2 62000_8000_M2 0.022
r 62000_8000_M2 62000_10000_M2 0.022
r 62000_10000_M2 62000_12000_M2 0.022
r 62000_12000_M2 62000_14000_M2 0.022
r 62000_14000_M2 62000_16000_M2 0.022
r 62000_16000_M2 62000_18000_M2 0.022
r 62000_18000_M2 62000_20000_M2 0.022
r 62000_20000_M2 62000_22000_M2 0.022
r 62000_22000_M2 62000_24000_M2 0.022
r 62000_24000_M2 62000_26000_M2 0.022
r 62000_26000_M2 62000_28000_M2 0.022
r 62000_28000_M2 62000_30000_M2 0.022
r 62000_30000_M2 62000_32000_M2 0.022
r 62000_32000_M2 62000_34000_M2 0.022
r 62000_34000_M2 62000_36000_M2 0.022
r 62000_36000_M2 62000_38000_M2 0.022
r 62000_38000_M2 62000_40000_M2 0.022
r 62000_40000_M2 62000_42000_M2 0.022
r 62000_42000_M2 62000_44000_M2 0.022
r 62000_44000_M2 62000_46000_M2 0.022
r 62000_46000_M2 62000_48000_M2 0.022
r 62000_48000_M2 62000_50000_M2 0.022
r 62000_50000_M2 62000_52000_M2 0.022
r 62000_52000_M2 62000_54000_M2 0.022
r 62000_54000_M2 62000_56000_M2 0.022
r 62000_56000_M2 62000_58000_M2 0.022
r 62000_58000_M2 62000_60000_M2 0.022
r 62000_60000_M2 62000_62000_M2 0.022
r 62000_62000_M2 62000_64000_M2 0.022
r 62000_64000_M2 62000_66000_M2 0.022
r 62000_66000_M2 62000_68000_M2 0.022
r 62000_68000_M2 62000_70000_M2 0.022
r 62000_70000_M2 62000_72000_M2 0.022
r 62000_72000_M2 62000_74000_M2 0.022
r 62000_74000_M2 62000_76000_M2 0.022
r 62000_76000_M2 62000_78000_M2 0.022
r 62000_78000_M2 62000_80000_M2 0.022
r 62000_80000_M2 62000_82000_M2 0.022
r 62000_82000_M2 62000_84000_M2 0.022
r 62000_84000_M2 62000_86000_M2 0.022
r 62000_86000_M2 62000_88000_M2 0.022
r 62000_88000_M2 62000_90000_M2 0.022
r 62000_90000_M2 62000_92000_M2 0.022
r 62000_92000_M2 62000_94000_M2 0.022
r 62000_94000_M2 62000_96000_M2 0.022
r 62000_96000_M2 62000_98000_M2 0.022
r 62000_98000_M2 62000_100000_M2 0.022
r 64000_2000_M2 64000_4000_M2 0.022
r 64000_4000_M2 64000_6000_M2 0.022
r 64000_6000_M2 64000_8000_M2 0.022
r 64000_8000_M2 64000_10000_M2 0.022
r 64000_10000_M2 64000_12000_M2 0.022
r 64000_12000_M2 64000_14000_M2 0.022
r 64000_14000_M2 64000_16000_M2 0.022
r 64000_16000_M2 64000_18000_M2 0.022
r 64000_18000_M2 64000_20000_M2 0.022
r 64000_20000_M2 64000_22000_M2 0.022
r 64000_22000_M2 64000_24000_M2 0.022
r 64000_24000_M2 64000_26000_M2 0.022
r 64000_26000_M2 64000_28000_M2 0.022
r 64000_28000_M2 64000_30000_M2 0.022
r 64000_30000_M2 64000_32000_M2 0.022
r 64000_32000_M2 64000_34000_M2 0.022
r 64000_34000_M2 64000_36000_M2 0.022
r 64000_36000_M2 64000_38000_M2 0.022
r 64000_38000_M2 64000_40000_M2 0.022
r 64000_40000_M2 64000_42000_M2 0.022
r 64000_42000_M2 64000_44000_M2 0.022
r 64000_44000_M2 64000_46000_M2 0.022
r 64000_46000_M2 64000_48000_M2 0.022
r 64000_48000_M2 64000_50000_M2 0.022
r 64000_50000_M2 64000_52000_M2 0.022
r 64000_52000_M2 64000_54000_M2 0.022
r 64000_54000_M2 64000_56000_M2 0.022
r 64000_56000_M2 64000_58000_M2 0.022
r 64000_58000_M2 64000_60000_M2 0.022
r 64000_60000_M2 64000_62000_M2 0.022
r 64000_62000_M2 64000_64000_M2 0.022
r 64000_64000_M2 64000_66000_M2 0.022
r 64000_66000_M2 64000_68000_M2 0.022
r 64000_68000_M2 64000_70000_M2 0.022
r 64000_70000_M2 64000_72000_M2 0.022
r 64000_72000_M2 64000_74000_M2 0.022
r 64000_74000_M2 64000_76000_M2 0.022
r 64000_76000_M2 64000_78000_M2 0.022
r 64000_78000_M2 64000_80000_M2 0.022
r 64000_80000_M2 64000_82000_M2 0.022
r 64000_82000_M2 64000_84000_M2 0.022
r 64000_84000_M2 64000_86000_M2 0.022
r 64000_86000_M2 64000_88000_M2 0.022
r 64000_88000_M2 64000_90000_M2 0.022
r 64000_90000_M2 64000_92000_M2 0.022
r 64000_92000_M2 64000_94000_M2 0.022
r 64000_94000_M2 64000_96000_M2 0.022
r 64000_96000_M2 64000_98000_M2 0.022
r 64000_98000_M2 64000_100000_M2 0.022
r 66000_2000_M2 66000_4000_M2 0.022
r 66000_4000_M2 66000_6000_M2 0.022
r 66000_6000_M2 66000_8000_M2 0.022
r 66000_8000_M2 66000_10000_M2 0.022
r 66000_10000_M2 66000_12000_M2 0.022
r 66000_12000_M2 66000_14000_M2 0.022
r 66000_14000_M2 66000_16000_M2 0.022
r 66000_16000_M2 66000_18000_M2 0.022
r 66000_18000_M2 66000_20000_M2 0.022
r 66000_20000_M2 66000_22000_M2 0.022
r 66000_22000_M2 66000_24000_M2 0.022
r 66000_24000_M2 66000_26000_M2 0.022
r 66000_26000_M2 66000_28000_M2 0.022
r 66000_28000_M2 66000_30000_M2 0.022
r 66000_30000_M2 66000_32000_M2 0.022
r 66000_32000_M2 66000_34000_M2 0.022
r 66000_34000_M2 66000_36000_M2 0.022
r 66000_36000_M2 66000_38000_M2 0.022
r 66000_38000_M2 66000_40000_M2 0.022
r 66000_40000_M2 66000_42000_M2 0.022
r 66000_42000_M2 66000_44000_M2 0.022
r 66000_44000_M2 66000_46000_M2 0.022
r 66000_46000_M2 66000_48000_M2 0.022
r 66000_48000_M2 66000_50000_M2 0.022
r 66000_50000_M2 66000_52000_M2 0.022
r 66000_52000_M2 66000_54000_M2 0.022
r 66000_54000_M2 66000_56000_M2 0.022
r 66000_56000_M2 66000_58000_M2 0.022
r 66000_58000_M2 66000_60000_M2 0.022
r 66000_60000_M2 66000_62000_M2 0.022
r 66000_62000_M2 66000_64000_M2 0.022
r 66000_64000_M2 66000_66000_M2 0.022
r 66000_66000_M2 66000_68000_M2 0.022
r 66000_68000_M2 66000_70000_M2 0.022
r 66000_70000_M2 66000_72000_M2 0.022
r 66000_72000_M2 66000_74000_M2 0.022
r 66000_74000_M2 66000_76000_M2 0.022
r 66000_76000_M2 66000_78000_M2 0.022
r 66000_78000_M2 66000_80000_M2 0.022
r 66000_80000_M2 66000_82000_M2 0.022
r 66000_82000_M2 66000_84000_M2 0.022
r 66000_84000_M2 66000_86000_M2 0.022
r 66000_86000_M2 66000_88000_M2 0.022
r 66000_88000_M2 66000_90000_M2 0.022
r 66000_90000_M2 66000_92000_M2 0.022
r 66000_92000_M2 66000_94000_M2 0.022
r 66000_94000_M2 66000_96000_M2 0.022
r 66000_96000_M2 66000_98000_M2 0.022
r 66000_98000_M2 66000_100000_M2 0.022
r 68000_2000_M2 68000_4000_M2 0.022
r 68000_4000_M2 68000_6000_M2 0.022
r 68000_6000_M2 68000_8000_M2 0.022
r 68000_8000_M2 68000_10000_M2 0.022
r 68000_10000_M2 68000_12000_M2 0.022
r 68000_12000_M2 68000_14000_M2 0.022
r 68000_14000_M2 68000_16000_M2 0.022
r 68000_16000_M2 68000_18000_M2 0.022
r 68000_18000_M2 68000_20000_M2 0.022
r 68000_20000_M2 68000_22000_M2 0.022
r 68000_22000_M2 68000_24000_M2 0.022
r 68000_24000_M2 68000_26000_M2 0.022
r 68000_26000_M2 68000_28000_M2 0.022
r 68000_28000_M2 68000_30000_M2 0.022
r 68000_30000_M2 68000_32000_M2 0.022
r 68000_32000_M2 68000_34000_M2 0.022
r 68000_34000_M2 68000_36000_M2 0.022
r 68000_36000_M2 68000_38000_M2 0.022
r 68000_38000_M2 68000_40000_M2 0.022
r 68000_40000_M2 68000_42000_M2 0.022
r 68000_42000_M2 68000_44000_M2 0.022
r 68000_44000_M2 68000_46000_M2 0.022
r 68000_46000_M2 68000_48000_M2 0.022
r 68000_48000_M2 68000_50000_M2 0.022
r 68000_50000_M2 68000_52000_M2 0.022
r 68000_52000_M2 68000_54000_M2 0.022
r 68000_54000_M2 68000_56000_M2 0.022
r 68000_56000_M2 68000_58000_M2 0.022
r 68000_58000_M2 68000_60000_M2 0.022
r 68000_60000_M2 68000_62000_M2 0.022
r 68000_62000_M2 68000_64000_M2 0.022
r 68000_64000_M2 68000_66000_M2 0.022
r 68000_66000_M2 68000_68000_M2 0.022
r 68000_68000_M2 68000_70000_M2 0.022
r 68000_70000_M2 68000_72000_M2 0.022
r 68000_72000_M2 68000_74000_M2 0.022
r 68000_74000_M2 68000_76000_M2 0.022
r 68000_76000_M2 68000_78000_M2 0.022
r 68000_78000_M2 68000_80000_M2 0.022
r 68000_80000_M2 68000_82000_M2 0.022
r 68000_82000_M2 68000_84000_M2 0.022
r 68000_84000_M2 68000_86000_M2 0.022
r 68000_86000_M2 68000_88000_M2 0.022
r 68000_88000_M2 68000_90000_M2 0.022
r 68000_90000_M2 68000_92000_M2 0.022
r 68000_92000_M2 68000_94000_M2 0.022
r 68000_94000_M2 68000_96000_M2 0.022
r 68000_96000_M2 68000_98000_M2 0.022
r 68000_98000_M2 68000_100000_M2 0.022
r 70000_2000_M2 70000_4000_M2 0.022
r 70000_4000_M2 70000_6000_M2 0.022
r 70000_6000_M2 70000_8000_M2 0.022
r 70000_8000_M2 70000_10000_M2 0.022
r 70000_10000_M2 70000_12000_M2 0.022
r 70000_12000_M2 70000_14000_M2 0.022
r 70000_14000_M2 70000_16000_M2 0.022
r 70000_16000_M2 70000_18000_M2 0.022
r 70000_18000_M2 70000_20000_M2 0.022
r 70000_20000_M2 70000_22000_M2 0.022
r 70000_22000_M2 70000_24000_M2 0.022
r 70000_24000_M2 70000_26000_M2 0.022
r 70000_26000_M2 70000_28000_M2 0.022
r 70000_28000_M2 70000_30000_M2 0.022
r 70000_30000_M2 70000_32000_M2 0.022
r 70000_32000_M2 70000_34000_M2 0.022
r 70000_34000_M2 70000_36000_M2 0.022
r 70000_36000_M2 70000_38000_M2 0.022
r 70000_38000_M2 70000_40000_M2 0.022
r 70000_40000_M2 70000_42000_M2 0.022
r 70000_42000_M2 70000_44000_M2 0.022
r 70000_44000_M2 70000_46000_M2 0.022
r 70000_46000_M2 70000_48000_M2 0.022
r 70000_48000_M2 70000_50000_M2 0.022
r 70000_50000_M2 70000_52000_M2 0.022
r 70000_52000_M2 70000_54000_M2 0.022
r 70000_54000_M2 70000_56000_M2 0.022
r 70000_56000_M2 70000_58000_M2 0.022
r 70000_58000_M2 70000_60000_M2 0.022
r 70000_60000_M2 70000_62000_M2 0.022
r 70000_62000_M2 70000_64000_M2 0.022
r 70000_64000_M2 70000_66000_M2 0.022
r 70000_66000_M2 70000_68000_M2 0.022
r 70000_68000_M2 70000_70000_M2 0.022
r 70000_70000_M2 70000_72000_M2 0.022
r 70000_72000_M2 70000_74000_M2 0.022
r 70000_74000_M2 70000_76000_M2 0.022
r 70000_76000_M2 70000_78000_M2 0.022
r 70000_78000_M2 70000_80000_M2 0.022
r 70000_80000_M2 70000_82000_M2 0.022
r 70000_82000_M2 70000_84000_M2 0.022
r 70000_84000_M2 70000_86000_M2 0.022
r 70000_86000_M2 70000_88000_M2 0.022
r 70000_88000_M2 70000_90000_M2 0.022
r 70000_90000_M2 70000_92000_M2 0.022
r 70000_92000_M2 70000_94000_M2 0.022
r 70000_94000_M2 70000_96000_M2 0.022
r 70000_96000_M2 70000_98000_M2 0.022
r 70000_98000_M2 70000_100000_M2 0.022
r 72000_2000_M2 72000_4000_M2 0.022
r 72000_4000_M2 72000_6000_M2 0.022
r 72000_6000_M2 72000_8000_M2 0.022
r 72000_8000_M2 72000_10000_M2 0.022
r 72000_10000_M2 72000_12000_M2 0.022
r 72000_12000_M2 72000_14000_M2 0.022
r 72000_14000_M2 72000_16000_M2 0.022
r 72000_16000_M2 72000_18000_M2 0.022
r 72000_18000_M2 72000_20000_M2 0.022
r 72000_20000_M2 72000_22000_M2 0.022
r 72000_22000_M2 72000_24000_M2 0.022
r 72000_24000_M2 72000_26000_M2 0.022
r 72000_26000_M2 72000_28000_M2 0.022
r 72000_28000_M2 72000_30000_M2 0.022
r 72000_30000_M2 72000_32000_M2 0.022
r 72000_32000_M2 72000_34000_M2 0.022
r 72000_34000_M2 72000_36000_M2 0.022
r 72000_36000_M2 72000_38000_M2 0.022
r 72000_38000_M2 72000_40000_M2 0.022
r 72000_40000_M2 72000_42000_M2 0.022
r 72000_42000_M2 72000_44000_M2 0.022
r 72000_44000_M2 72000_46000_M2 0.022
r 72000_46000_M2 72000_48000_M2 0.022
r 72000_48000_M2 72000_50000_M2 0.022
r 72000_50000_M2 72000_52000_M2 0.022
r 72000_52000_M2 72000_54000_M2 0.022
r 72000_54000_M2 72000_56000_M2 0.022
r 72000_56000_M2 72000_58000_M2 0.022
r 72000_58000_M2 72000_60000_M2 0.022
r 72000_60000_M2 72000_62000_M2 0.022
r 72000_62000_M2 72000_64000_M2 0.022
r 72000_64000_M2 72000_66000_M2 0.022
r 72000_66000_M2 72000_68000_M2 0.022
r 72000_68000_M2 72000_70000_M2 0.022
r 72000_70000_M2 72000_72000_M2 0.022
r 72000_72000_M2 72000_74000_M2 0.022
r 72000_74000_M2 72000_76000_M2 0.022
r 72000_76000_M2 72000_78000_M2 0.022
r 72000_78000_M2 72000_80000_M2 0.022
r 72000_80000_M2 72000_82000_M2 0.022
r 72000_82000_M2 72000_84000_M2 0.022
r 72000_84000_M2 72000_86000_M2 0.022
r 72000_86000_M2 72000_88000_M2 0.022
r 72000_88000_M2 72000_90000_M2 0.022
r 72000_90000_M2 72000_92000_M2 0.022
r 72000_92000_M2 72000_94000_M2 0.022
r 72000_94000_M2 72000_96000_M2 0.022
r 72000_96000_M2 72000_98000_M2 0.022
r 72000_98000_M2 72000_100000_M2 0.022
r 74000_2000_M2 74000_4000_M2 0.022
r 74000_4000_M2 74000_6000_M2 0.022
r 74000_6000_M2 74000_8000_M2 0.022
r 74000_8000_M2 74000_10000_M2 0.022
r 74000_10000_M2 74000_12000_M2 0.022
r 74000_12000_M2 74000_14000_M2 0.022
r 74000_14000_M2 74000_16000_M2 0.022
r 74000_16000_M2 74000_18000_M2 0.022
r 74000_18000_M2 74000_20000_M2 0.022
r 74000_20000_M2 74000_22000_M2 0.022
r 74000_22000_M2 74000_24000_M2 0.022
r 74000_24000_M2 74000_26000_M2 0.022
r 74000_26000_M2 74000_28000_M2 0.022
r 74000_28000_M2 74000_30000_M2 0.022
r 74000_30000_M2 74000_32000_M2 0.022
r 74000_32000_M2 74000_34000_M2 0.022
r 74000_34000_M2 74000_36000_M2 0.022
r 74000_36000_M2 74000_38000_M2 0.022
r 74000_38000_M2 74000_40000_M2 0.022
r 74000_40000_M2 74000_42000_M2 0.022
r 74000_42000_M2 74000_44000_M2 0.022
r 74000_44000_M2 74000_46000_M2 0.022
r 74000_46000_M2 74000_48000_M2 0.022
r 74000_48000_M2 74000_50000_M2 0.022
r 74000_50000_M2 74000_52000_M2 0.022
r 74000_52000_M2 74000_54000_M2 0.022
r 74000_54000_M2 74000_56000_M2 0.022
r 74000_56000_M2 74000_58000_M2 0.022
r 74000_58000_M2 74000_60000_M2 0.022
r 74000_60000_M2 74000_62000_M2 0.022
r 74000_62000_M2 74000_64000_M2 0.022
r 74000_64000_M2 74000_66000_M2 0.022
r 74000_66000_M2 74000_68000_M2 0.022
r 74000_68000_M2 74000_70000_M2 0.022
r 74000_70000_M2 74000_72000_M2 0.022
r 74000_72000_M2 74000_74000_M2 0.022
r 74000_74000_M2 74000_76000_M2 0.022
r 74000_76000_M2 74000_78000_M2 0.022
r 74000_78000_M2 74000_80000_M2 0.022
r 74000_80000_M2 74000_82000_M2 0.022
r 74000_82000_M2 74000_84000_M2 0.022
r 74000_84000_M2 74000_86000_M2 0.022
r 74000_86000_M2 74000_88000_M2 0.022
r 74000_88000_M2 74000_90000_M2 0.022
r 74000_90000_M2 74000_92000_M2 0.022
r 74000_92000_M2 74000_94000_M2 0.022
r 74000_94000_M2 74000_96000_M2 0.022
r 74000_96000_M2 74000_98000_M2 0.022
r 74000_98000_M2 74000_100000_M2 0.022
r 76000_2000_M2 76000_4000_M2 0.022
r 76000_4000_M2 76000_6000_M2 0.022
r 76000_6000_M2 76000_8000_M2 0.022
r 76000_8000_M2 76000_10000_M2 0.022
r 76000_10000_M2 76000_12000_M2 0.022
r 76000_12000_M2 76000_14000_M2 0.022
r 76000_14000_M2 76000_16000_M2 0.022
r 76000_16000_M2 76000_18000_M2 0.022
r 76000_18000_M2 76000_20000_M2 0.022
r 76000_20000_M2 76000_22000_M2 0.022
r 76000_22000_M2 76000_24000_M2 0.022
r 76000_24000_M2 76000_26000_M2 0.022
r 76000_26000_M2 76000_28000_M2 0.022
r 76000_28000_M2 76000_30000_M2 0.022
r 76000_30000_M2 76000_32000_M2 0.022
r 76000_32000_M2 76000_34000_M2 0.022
r 76000_34000_M2 76000_36000_M2 0.022
r 76000_36000_M2 76000_38000_M2 0.022
r 76000_38000_M2 76000_40000_M2 0.022
r 76000_40000_M2 76000_42000_M2 0.022
r 76000_42000_M2 76000_44000_M2 0.022
r 76000_44000_M2 76000_46000_M2 0.022
r 76000_46000_M2 76000_48000_M2 0.022
r 76000_48000_M2 76000_50000_M2 0.022
r 76000_50000_M2 76000_52000_M2 0.022
r 76000_52000_M2 76000_54000_M2 0.022
r 76000_54000_M2 76000_56000_M2 0.022
r 76000_56000_M2 76000_58000_M2 0.022
r 76000_58000_M2 76000_60000_M2 0.022
r 76000_60000_M2 76000_62000_M2 0.022
r 76000_62000_M2 76000_64000_M2 0.022
r 76000_64000_M2 76000_66000_M2 0.022
r 76000_66000_M2 76000_68000_M2 0.022
r 76000_68000_M2 76000_70000_M2 0.022
r 76000_70000_M2 76000_72000_M2 0.022
r 76000_72000_M2 76000_74000_M2 0.022
r 76000_74000_M2 76000_76000_M2 0.022
r 76000_76000_M2 76000_78000_M2 0.022
r 76000_78000_M2 76000_80000_M2 0.022
r 76000_80000_M2 76000_82000_M2 0.022
r 76000_82000_M2 76000_84000_M2 0.022
r 76000_84000_M2 76000_86000_M2 0.022
r 76000_86000_M2 76000_88000_M2 0.022
r 76000_88000_M2 76000_90000_M2 0.022
r 76000_90000_M2 76000_92000_M2 0.022
r 76000_92000_M2 76000_94000_M2 0.022
r 76000_94000_M2 76000_96000_M2 0.022
r 76000_96000_M2 76000_98000_M2 0.022
r 76000_98000_M2 76000_100000_M2 0.022
r 78000_2000_M2 78000_4000_M2 0.022
r 78000_4000_M2 78000_6000_M2 0.022
r 78000_6000_M2 78000_8000_M2 0.022
r 78000_8000_M2 78000_10000_M2 0.022
r 78000_10000_M2 78000_12000_M2 0.022
r 78000_12000_M2 78000_14000_M2 0.022
r 78000_14000_M2 78000_16000_M2 0.022
r 78000_16000_M2 78000_18000_M2 0.022
r 78000_18000_M2 78000_20000_M2 0.022
r 78000_20000_M2 78000_22000_M2 0.022
r 78000_22000_M2 78000_24000_M2 0.022
r 78000_24000_M2 78000_26000_M2 0.022
r 78000_26000_M2 78000_28000_M2 0.022
r 78000_28000_M2 78000_30000_M2 0.022
r 78000_30000_M2 78000_32000_M2 0.022
r 78000_32000_M2 78000_34000_M2 0.022
r 78000_34000_M2 78000_36000_M2 0.022
r 78000_36000_M2 78000_38000_M2 0.022
r 78000_38000_M2 78000_40000_M2 0.022
r 78000_40000_M2 78000_42000_M2 0.022
r 78000_42000_M2 78000_44000_M2 0.022
r 78000_44000_M2 78000_46000_M2 0.022
r 78000_46000_M2 78000_48000_M2 0.022
r 78000_48000_M2 78000_50000_M2 0.022
r 78000_50000_M2 78000_52000_M2 0.022
r 78000_52000_M2 78000_54000_M2 0.022
r 78000_54000_M2 78000_56000_M2 0.022
r 78000_56000_M2 78000_58000_M2 0.022
r 78000_58000_M2 78000_60000_M2 0.022
r 78000_60000_M2 78000_62000_M2 0.022
r 78000_62000_M2 78000_64000_M2 0.022
r 78000_64000_M2 78000_66000_M2 0.022
r 78000_66000_M2 78000_68000_M2 0.022
r 78000_68000_M2 78000_70000_M2 0.022
r 78000_70000_M2 78000_72000_M2 0.022
r 78000_72000_M2 78000_74000_M2 0.022
r 78000_74000_M2 78000_76000_M2 0.022
r 78000_76000_M2 78000_78000_M2 0.022
r 78000_78000_M2 78000_80000_M2 0.022
r 78000_80000_M2 78000_82000_M2 0.022
r 78000_82000_M2 78000_84000_M2 0.022
r 78000_84000_M2 78000_86000_M2 0.022
r 78000_86000_M2 78000_88000_M2 0.022
r 78000_88000_M2 78000_90000_M2 0.022
r 78000_90000_M2 78000_92000_M2 0.022
r 78000_92000_M2 78000_94000_M2 0.022
r 78000_94000_M2 78000_96000_M2 0.022
r 78000_96000_M2 78000_98000_M2 0.022
r 78000_98000_M2 78000_100000_M2 0.022
r 80000_2000_M2 80000_4000_M2 0.022
r 80000_4000_M2 80000_6000_M2 0.022
r 80000_6000_M2 80000_8000_M2 0.022
r 80000_8000_M2 80000_10000_M2 0.022
r 80000_10000_M2 80000_12000_M2 0.022
r 80000_12000_M2 80000_14000_M2 0.022
r 80000_14000_M2 80000_16000_M2 0.022
r 80000_16000_M2 80000_18000_M2 0.022
r 80000_18000_M2 80000_20000_M2 0.022
r 80000_20000_M2 80000_22000_M2 0.022
r 80000_22000_M2 80000_24000_M2 0.022
r 80000_24000_M2 80000_26000_M2 0.022
r 80000_26000_M2 80000_28000_M2 0.022
r 80000_28000_M2 80000_30000_M2 0.022
r 80000_30000_M2 80000_32000_M2 0.022
r 80000_32000_M2 80000_34000_M2 0.022
r 80000_34000_M2 80000_36000_M2 0.022
r 80000_36000_M2 80000_38000_M2 0.022
r 80000_38000_M2 80000_40000_M2 0.022
r 80000_40000_M2 80000_42000_M2 0.022
r 80000_42000_M2 80000_44000_M2 0.022
r 80000_44000_M2 80000_46000_M2 0.022
r 80000_46000_M2 80000_48000_M2 0.022
r 80000_48000_M2 80000_50000_M2 0.022
r 80000_50000_M2 80000_52000_M2 0.022
r 80000_52000_M2 80000_54000_M2 0.022
r 80000_54000_M2 80000_56000_M2 0.022
r 80000_56000_M2 80000_58000_M2 0.022
r 80000_58000_M2 80000_60000_M2 0.022
r 80000_60000_M2 80000_62000_M2 0.022
r 80000_62000_M2 80000_64000_M2 0.022
r 80000_64000_M2 80000_66000_M2 0.022
r 80000_66000_M2 80000_68000_M2 0.022
r 80000_68000_M2 80000_70000_M2 0.022
r 80000_70000_M2 80000_72000_M2 0.022
r 80000_72000_M2 80000_74000_M2 0.022
r 80000_74000_M2 80000_76000_M2 0.022
r 80000_76000_M2 80000_78000_M2 0.022
r 80000_78000_M2 80000_80000_M2 0.022
r 80000_80000_M2 80000_82000_M2 0.022
r 80000_82000_M2 80000_84000_M2 0.022
r 80000_84000_M2 80000_86000_M2 0.022
r 80000_86000_M2 80000_88000_M2 0.022
r 80000_88000_M2 80000_90000_M2 0.022
r 80000_90000_M2 80000_92000_M2 0.022
r 80000_92000_M2 80000_94000_M2 0.022
r 80000_94000_M2 80000_96000_M2 0.022
r 80000_96000_M2 80000_98000_M2 0.022
r 80000_98000_M2 80000_100000_M2 0.022
r 82000_2000_M2 82000_4000_M2 0.022
r 82000_4000_M2 82000_6000_M2 0.022
r 82000_6000_M2 82000_8000_M2 0.022
r 82000_8000_M2 82000_10000_M2 0.022
r 82000_10000_M2 82000_12000_M2 0.022
r 82000_12000_M2 82000_14000_M2 0.022
r 82000_14000_M2 82000_16000_M2 0.022
r 82000_16000_M2 82000_18000_M2 0.022
r 82000_18000_M2 82000_20000_M2 0.022
r 82000_20000_M2 82000_22000_M2 0.022
r 82000_22000_M2 82000_24000_M2 0.022
r 82000_24000_M2 82000_26000_M2 0.022
r 82000_26000_M2 82000_28000_M2 0.022
r 82000_28000_M2 82000_30000_M2 0.022
r 82000_30000_M2 82000_32000_M2 0.022
r 82000_32000_M2 82000_34000_M2 0.022
r 82000_34000_M2 82000_36000_M2 0.022
r 82000_36000_M2 82000_38000_M2 0.022
r 82000_38000_M2 82000_40000_M2 0.022
r 82000_40000_M2 82000_42000_M2 0.022
r 82000_42000_M2 82000_44000_M2 0.022
r 82000_44000_M2 82000_46000_M2 0.022
r 82000_46000_M2 82000_48000_M2 0.022
r 82000_48000_M2 82000_50000_M2 0.022
r 82000_50000_M2 82000_52000_M2 0.022
r 82000_52000_M2 82000_54000_M2 0.022
r 82000_54000_M2 82000_56000_M2 0.022
r 82000_56000_M2 82000_58000_M2 0.022
r 82000_58000_M2 82000_60000_M2 0.022
r 82000_60000_M2 82000_62000_M2 0.022
r 82000_62000_M2 82000_64000_M2 0.022
r 82000_64000_M2 82000_66000_M2 0.022
r 82000_66000_M2 82000_68000_M2 0.022
r 82000_68000_M2 82000_70000_M2 0.022
r 82000_70000_M2 82000_72000_M2 0.022
r 82000_72000_M2 82000_74000_M2 0.022
r 82000_74000_M2 82000_76000_M2 0.022
r 82000_76000_M2 82000_78000_M2 0.022
r 82000_78000_M2 82000_80000_M2 0.022
r 82000_80000_M2 82000_82000_M2 0.022
r 82000_82000_M2 82000_84000_M2 0.022
r 82000_84000_M2 82000_86000_M2 0.022
r 82000_86000_M2 82000_88000_M2 0.022
r 82000_88000_M2 82000_90000_M2 0.022
r 82000_90000_M2 82000_92000_M2 0.022
r 82000_92000_M2 82000_94000_M2 0.022
r 82000_94000_M2 82000_96000_M2 0.022
r 82000_96000_M2 82000_98000_M2 0.022
r 82000_98000_M2 82000_100000_M2 0.022
r 84000_2000_M2 84000_4000_M2 0.022
r 84000_4000_M2 84000_6000_M2 0.022
r 84000_6000_M2 84000_8000_M2 0.022
r 84000_8000_M2 84000_10000_M2 0.022
r 84000_10000_M2 84000_12000_M2 0.022
r 84000_12000_M2 84000_14000_M2 0.022
r 84000_14000_M2 84000_16000_M2 0.022
r 84000_16000_M2 84000_18000_M2 0.022
r 84000_18000_M2 84000_20000_M2 0.022
r 84000_20000_M2 84000_22000_M2 0.022
r 84000_22000_M2 84000_24000_M2 0.022
r 84000_24000_M2 84000_26000_M2 0.022
r 84000_26000_M2 84000_28000_M2 0.022
r 84000_28000_M2 84000_30000_M2 0.022
r 84000_30000_M2 84000_32000_M2 0.022
r 84000_32000_M2 84000_34000_M2 0.022
r 84000_34000_M2 84000_36000_M2 0.022
r 84000_36000_M2 84000_38000_M2 0.022
r 84000_38000_M2 84000_40000_M2 0.022
r 84000_40000_M2 84000_42000_M2 0.022
r 84000_42000_M2 84000_44000_M2 0.022
r 84000_44000_M2 84000_46000_M2 0.022
r 84000_46000_M2 84000_48000_M2 0.022
r 84000_48000_M2 84000_50000_M2 0.022
r 84000_50000_M2 84000_52000_M2 0.022
r 84000_52000_M2 84000_54000_M2 0.022
r 84000_54000_M2 84000_56000_M2 0.022
r 84000_56000_M2 84000_58000_M2 0.022
r 84000_58000_M2 84000_60000_M2 0.022
r 84000_60000_M2 84000_62000_M2 0.022
r 84000_62000_M2 84000_64000_M2 0.022
r 84000_64000_M2 84000_66000_M2 0.022
r 84000_66000_M2 84000_68000_M2 0.022
r 84000_68000_M2 84000_70000_M2 0.022
r 84000_70000_M2 84000_72000_M2 0.022
r 84000_72000_M2 84000_74000_M2 0.022
r 84000_74000_M2 84000_76000_M2 0.022
r 84000_76000_M2 84000_78000_M2 0.022
r 84000_78000_M2 84000_80000_M2 0.022
r 84000_80000_M2 84000_82000_M2 0.022
r 84000_82000_M2 84000_84000_M2 0.022
r 84000_84000_M2 84000_86000_M2 0.022
r 84000_86000_M2 84000_88000_M2 0.022
r 84000_88000_M2 84000_90000_M2 0.022
r 84000_90000_M2 84000_92000_M2 0.022
r 84000_92000_M2 84000_94000_M2 0.022
r 84000_94000_M2 84000_96000_M2 0.022
r 84000_96000_M2 84000_98000_M2 0.022
r 84000_98000_M2 84000_100000_M2 0.022
r 86000_2000_M2 86000_4000_M2 0.022
r 86000_4000_M2 86000_6000_M2 0.022
r 86000_6000_M2 86000_8000_M2 0.022
r 86000_8000_M2 86000_10000_M2 0.022
r 86000_10000_M2 86000_12000_M2 0.022
r 86000_12000_M2 86000_14000_M2 0.022
r 86000_14000_M2 86000_16000_M2 0.022
r 86000_16000_M2 86000_18000_M2 0.022
r 86000_18000_M2 86000_20000_M2 0.022
r 86000_20000_M2 86000_22000_M2 0.022
r 86000_22000_M2 86000_24000_M2 0.022
r 86000_24000_M2 86000_26000_M2 0.022
r 86000_26000_M2 86000_28000_M2 0.022
r 86000_28000_M2 86000_30000_M2 0.022
r 86000_30000_M2 86000_32000_M2 0.022
r 86000_32000_M2 86000_34000_M2 0.022
r 86000_34000_M2 86000_36000_M2 0.022
r 86000_36000_M2 86000_38000_M2 0.022
r 86000_38000_M2 86000_40000_M2 0.022
r 86000_40000_M2 86000_42000_M2 0.022
r 86000_42000_M2 86000_44000_M2 0.022
r 86000_44000_M2 86000_46000_M2 0.022
r 86000_46000_M2 86000_48000_M2 0.022
r 86000_48000_M2 86000_50000_M2 0.022
r 86000_50000_M2 86000_52000_M2 0.022
r 86000_52000_M2 86000_54000_M2 0.022
r 86000_54000_M2 86000_56000_M2 0.022
r 86000_56000_M2 86000_58000_M2 0.022
r 86000_58000_M2 86000_60000_M2 0.022
r 86000_60000_M2 86000_62000_M2 0.022
r 86000_62000_M2 86000_64000_M2 0.022
r 86000_64000_M2 86000_66000_M2 0.022
r 86000_66000_M2 86000_68000_M2 0.022
r 86000_68000_M2 86000_70000_M2 0.022
r 86000_70000_M2 86000_72000_M2 0.022
r 86000_72000_M2 86000_74000_M2 0.022
r 86000_74000_M2 86000_76000_M2 0.022
r 86000_76000_M2 86000_78000_M2 0.022
r 86000_78000_M2 86000_80000_M2 0.022
r 86000_80000_M2 86000_82000_M2 0.022
r 86000_82000_M2 86000_84000_M2 0.022
r 86000_84000_M2 86000_86000_M2 0.022
r 86000_86000_M2 86000_88000_M2 0.022
r 86000_88000_M2 86000_90000_M2 0.022
r 86000_90000_M2 86000_92000_M2 0.022
r 86000_92000_M2 86000_94000_M2 0.022
r 86000_94000_M2 86000_96000_M2 0.022
r 86000_96000_M2 86000_98000_M2 0.022
r 86000_98000_M2 86000_100000_M2 0.022
r 88000_2000_M2 88000_4000_M2 0.022
r 88000_4000_M2 88000_6000_M2 0.022
r 88000_6000_M2 88000_8000_M2 0.022
r 88000_8000_M2 88000_10000_M2 0.022
r 88000_10000_M2 88000_12000_M2 0.022
r 88000_12000_M2 88000_14000_M2 0.022
r 88000_14000_M2 88000_16000_M2 0.022
r 88000_16000_M2 88000_18000_M2 0.022
r 88000_18000_M2 88000_20000_M2 0.022
r 88000_20000_M2 88000_22000_M2 0.022
r 88000_22000_M2 88000_24000_M2 0.022
r 88000_24000_M2 88000_26000_M2 0.022
r 88000_26000_M2 88000_28000_M2 0.022
r 88000_28000_M2 88000_30000_M2 0.022
r 88000_30000_M2 88000_32000_M2 0.022
r 88000_32000_M2 88000_34000_M2 0.022
r 88000_34000_M2 88000_36000_M2 0.022
r 88000_36000_M2 88000_38000_M2 0.022
r 88000_38000_M2 88000_40000_M2 0.022
r 88000_40000_M2 88000_42000_M2 0.022
r 88000_42000_M2 88000_44000_M2 0.022
r 88000_44000_M2 88000_46000_M2 0.022
r 88000_46000_M2 88000_48000_M2 0.022
r 88000_48000_M2 88000_50000_M2 0.022
r 88000_50000_M2 88000_52000_M2 0.022
r 88000_52000_M2 88000_54000_M2 0.022
r 88000_54000_M2 88000_56000_M2 0.022
r 88000_56000_M2 88000_58000_M2 0.022
r 88000_58000_M2 88000_60000_M2 0.022
r 88000_60000_M2 88000_62000_M2 0.022
r 88000_62000_M2 88000_64000_M2 0.022
r 88000_64000_M2 88000_66000_M2 0.022
r 88000_66000_M2 88000_68000_M2 0.022
r 88000_68000_M2 88000_70000_M2 0.022
r 88000_70000_M2 88000_72000_M2 0.022
r 88000_72000_M2 88000_74000_M2 0.022
r 88000_74000_M2 88000_76000_M2 0.022
r 88000_76000_M2 88000_78000_M2 0.022
r 88000_78000_M2 88000_80000_M2 0.022
r 88000_80000_M2 88000_82000_M2 0.022
r 88000_82000_M2 88000_84000_M2 0.022
r 88000_84000_M2 88000_86000_M2 0.022
r 88000_86000_M2 88000_88000_M2 0.022
r 88000_88000_M2 88000_90000_M2 0.022
r 88000_90000_M2 88000_92000_M2 0.022
r 88000_92000_M2 88000_94000_M2 0.022
r 88000_94000_M2 88000_96000_M2 0.022
r 88000_96000_M2 88000_98000_M2 0.022
r 88000_98000_M2 88000_100000_M2 0.022
r 90000_2000_M2 90000_4000_M2 0.022
r 90000_4000_M2 90000_6000_M2 0.022
r 90000_6000_M2 90000_8000_M2 0.022
r 90000_8000_M2 90000_10000_M2 0.022
r 90000_10000_M2 90000_12000_M2 0.022
r 90000_12000_M2 90000_14000_M2 0.022
r 90000_14000_M2 90000_16000_M2 0.022
r 90000_16000_M2 90000_18000_M2 0.022
r 90000_18000_M2 90000_20000_M2 0.022
r 90000_20000_M2 90000_22000_M2 0.022
r 90000_22000_M2 90000_24000_M2 0.022
r 90000_24000_M2 90000_26000_M2 0.022
r 90000_26000_M2 90000_28000_M2 0.022
r 90000_28000_M2 90000_30000_M2 0.022
r 90000_30000_M2 90000_32000_M2 0.022
r 90000_32000_M2 90000_34000_M2 0.022
r 90000_34000_M2 90000_36000_M2 0.022
r 90000_36000_M2 90000_38000_M2 0.022
r 90000_38000_M2 90000_40000_M2 0.022
r 90000_40000_M2 90000_42000_M2 0.022
r 90000_42000_M2 90000_44000_M2 0.022
r 90000_44000_M2 90000_46000_M2 0.022
r 90000_46000_M2 90000_48000_M2 0.022
r 90000_48000_M2 90000_50000_M2 0.022
r 90000_50000_M2 90000_52000_M2 0.022
r 90000_52000_M2 90000_54000_M2 0.022
r 90000_54000_M2 90000_56000_M2 0.022
r 90000_56000_M2 90000_58000_M2 0.022
r 90000_58000_M2 90000_60000_M2 0.022
r 90000_60000_M2 90000_62000_M2 0.022
r 90000_62000_M2 90000_64000_M2 0.022
r 90000_64000_M2 90000_66000_M2 0.022
r 90000_66000_M2 90000_68000_M2 0.022
r 90000_68000_M2 90000_70000_M2 0.022
r 90000_70000_M2 90000_72000_M2 0.022
r 90000_72000_M2 90000_74000_M2 0.022
r 90000_74000_M2 90000_76000_M2 0.022
r 90000_76000_M2 90000_78000_M2 0.022
r 90000_78000_M2 90000_80000_M2 0.022
r 90000_80000_M2 90000_82000_M2 0.022
r 90000_82000_M2 90000_84000_M2 0.022
r 90000_84000_M2 90000_86000_M2 0.022
r 90000_86000_M2 90000_88000_M2 0.022
r 90000_88000_M2 90000_90000_M2 0.022
r 90000_90000_M2 90000_92000_M2 0.022
r 90000_92000_M2 90000_94000_M2 0.022
r 90000_94000_M2 90000_96000_M2 0.022
r 90000_96000_M2 90000_98000_M2 0.022
r 90000_98000_M2 90000_100000_M2 0.022
r 92000_2000_M2 92000_4000_M2 0.022
r 92000_4000_M2 92000_6000_M2 0.022
r 92000_6000_M2 92000_8000_M2 0.022
r 92000_8000_M2 92000_10000_M2 0.022
r 92000_10000_M2 92000_12000_M2 0.022
r 92000_12000_M2 92000_14000_M2 0.022
r 92000_14000_M2 92000_16000_M2 0.022
r 92000_16000_M2 92000_18000_M2 0.022
r 92000_18000_M2 92000_20000_M2 0.022
r 92000_20000_M2 92000_22000_M2 0.022
r 92000_22000_M2 92000_24000_M2 0.022
r 92000_24000_M2 92000_26000_M2 0.022
r 92000_26000_M2 92000_28000_M2 0.022
r 92000_28000_M2 92000_30000_M2 0.022
r 92000_30000_M2 92000_32000_M2 0.022
r 92000_32000_M2 92000_34000_M2 0.022
r 92000_34000_M2 92000_36000_M2 0.022
r 92000_36000_M2 92000_38000_M2 0.022
r 92000_38000_M2 92000_40000_M2 0.022
r 92000_40000_M2 92000_42000_M2 0.022
r 92000_42000_M2 92000_44000_M2 0.022
r 92000_44000_M2 92000_46000_M2 0.022
r 92000_46000_M2 92000_48000_M2 0.022
r 92000_48000_M2 92000_50000_M2 0.022
r 92000_50000_M2 92000_52000_M2 0.022
r 92000_52000_M2 92000_54000_M2 0.022
r 92000_54000_M2 92000_56000_M2 0.022
r 92000_56000_M2 92000_58000_M2 0.022
r 92000_58000_M2 92000_60000_M2 0.022
r 92000_60000_M2 92000_62000_M2 0.022
r 92000_62000_M2 92000_64000_M2 0.022
r 92000_64000_M2 92000_66000_M2 0.022
r 92000_66000_M2 92000_68000_M2 0.022
r 92000_68000_M2 92000_70000_M2 0.022
r 92000_70000_M2 92000_72000_M2 0.022
r 92000_72000_M2 92000_74000_M2 0.022
r 92000_74000_M2 92000_76000_M2 0.022
r 92000_76000_M2 92000_78000_M2 0.022
r 92000_78000_M2 92000_80000_M2 0.022
r 92000_80000_M2 92000_82000_M2 0.022
r 92000_82000_M2 92000_84000_M2 0.022
r 92000_84000_M2 92000_86000_M2 0.022
r 92000_86000_M2 92000_88000_M2 0.022
r 92000_88000_M2 92000_90000_M2 0.022
r 92000_90000_M2 92000_92000_M2 0.022
r 92000_92000_M2 92000_94000_M2 0.022
r 92000_94000_M2 92000_96000_M2 0.022
r 92000_96000_M2 92000_98000_M2 0.022
r 92000_98000_M2 92000_100000_M2 0.022
r 94000_2000_M2 94000_4000_M2 0.022
r 94000_4000_M2 94000_6000_M2 0.022
r 94000_6000_M2 94000_8000_M2 0.022
r 94000_8000_M2 94000_10000_M2 0.022
r 94000_10000_M2 94000_12000_M2 0.022
r 94000_12000_M2 94000_14000_M2 0.022
r 94000_14000_M2 94000_16000_M2 0.022
r 94000_16000_M2 94000_18000_M2 0.022
r 94000_18000_M2 94000_20000_M2 0.022
r 94000_20000_M2 94000_22000_M2 0.022
r 94000_22000_M2 94000_24000_M2 0.022
r 94000_24000_M2 94000_26000_M2 0.022
r 94000_26000_M2 94000_28000_M2 0.022
r 94000_28000_M2 94000_30000_M2 0.022
r 94000_30000_M2 94000_32000_M2 0.022
r 94000_32000_M2 94000_34000_M2 0.022
r 94000_34000_M2 94000_36000_M2 0.022
r 94000_36000_M2 94000_38000_M2 0.022
r 94000_38000_M2 94000_40000_M2 0.022
r 94000_40000_M2 94000_42000_M2 0.022
r 94000_42000_M2 94000_44000_M2 0.022
r 94000_44000_M2 94000_46000_M2 0.022
r 94000_46000_M2 94000_48000_M2 0.022
r 94000_48000_M2 94000_50000_M2 0.022
r 94000_50000_M2 94000_52000_M2 0.022
r 94000_52000_M2 94000_54000_M2 0.022
r 94000_54000_M2 94000_56000_M2 0.022
r 94000_56000_M2 94000_58000_M2 0.022
r 94000_58000_M2 94000_60000_M2 0.022
r 94000_60000_M2 94000_62000_M2 0.022
r 94000_62000_M2 94000_64000_M2 0.022
r 94000_64000_M2 94000_66000_M2 0.022
r 94000_66000_M2 94000_68000_M2 0.022
r 94000_68000_M2 94000_70000_M2 0.022
r 94000_70000_M2 94000_72000_M2 0.022
r 94000_72000_M2 94000_74000_M2 0.022
r 94000_74000_M2 94000_76000_M2 0.022
r 94000_76000_M2 94000_78000_M2 0.022
r 94000_78000_M2 94000_80000_M2 0.022
r 94000_80000_M2 94000_82000_M2 0.022
r 94000_82000_M2 94000_84000_M2 0.022
r 94000_84000_M2 94000_86000_M2 0.022
r 94000_86000_M2 94000_88000_M2 0.022
r 94000_88000_M2 94000_90000_M2 0.022
r 94000_90000_M2 94000_92000_M2 0.022
r 94000_92000_M2 94000_94000_M2 0.022
r 94000_94000_M2 94000_96000_M2 0.022
r 94000_96000_M2 94000_98000_M2 0.022
r 94000_98000_M2 94000_100000_M2 0.022
r 96000_2000_M2 96000_4000_M2 0.022
r 96000_4000_M2 96000_6000_M2 0.022
r 96000_6000_M2 96000_8000_M2 0.022
r 96000_8000_M2 96000_10000_M2 0.022
r 96000_10000_M2 96000_12000_M2 0.022
r 96000_12000_M2 96000_14000_M2 0.022
r 96000_14000_M2 96000_16000_M2 0.022
r 96000_16000_M2 96000_18000_M2 0.022
r 96000_18000_M2 96000_20000_M2 0.022
r 96000_20000_M2 96000_22000_M2 0.022
r 96000_22000_M2 96000_24000_M2 0.022
r 96000_24000_M2 96000_26000_M2 0.022
r 96000_26000_M2 96000_28000_M2 0.022
r 96000_28000_M2 96000_30000_M2 0.022
r 96000_30000_M2 96000_32000_M2 0.022
r 96000_32000_M2 96000_34000_M2 0.022
r 96000_34000_M2 96000_36000_M2 0.022
r 96000_36000_M2 96000_38000_M2 0.022
r 96000_38000_M2 96000_40000_M2 0.022
r 96000_40000_M2 96000_42000_M2 0.022
r 96000_42000_M2 96000_44000_M2 0.022
r 96000_44000_M2 96000_46000_M2 0.022
r 96000_46000_M2 96000_48000_M2 0.022
r 96000_48000_M2 96000_50000_M2 0.022
r 96000_50000_M2 96000_52000_M2 0.022
r 96000_52000_M2 96000_54000_M2 0.022
r 96000_54000_M2 96000_56000_M2 0.022
r 96000_56000_M2 96000_58000_M2 0.022
r 96000_58000_M2 96000_60000_M2 0.022
r 96000_60000_M2 96000_62000_M2 0.022
r 96000_62000_M2 96000_64000_M2 0.022
r 96000_64000_M2 96000_66000_M2 0.022
r 96000_66000_M2 96000_68000_M2 0.022
r 96000_68000_M2 96000_70000_M2 0.022
r 96000_70000_M2 96000_72000_M2 0.022
r 96000_72000_M2 96000_74000_M2 0.022
r 96000_74000_M2 96000_76000_M2 0.022
r 96000_76000_M2 96000_78000_M2 0.022
r 96000_78000_M2 96000_80000_M2 0.022
r 96000_80000_M2 96000_82000_M2 0.022
r 96000_82000_M2 96000_84000_M2 0.022
r 96000_84000_M2 96000_86000_M2 0.022
r 96000_86000_M2 96000_88000_M2 0.022
r 96000_88000_M2 96000_90000_M2 0.022
r 96000_90000_M2 96000_92000_M2 0.022
r 96000_92000_M2 96000_94000_M2 0.022
r 96000_94000_M2 96000_96000_M2 0.022
r 96000_96000_M2 96000_98000_M2 0.022
r 96000_98000_M2 96000_100000_M2 0.022
r 98000_2000_M2 98000_4000_M2 0.022
r 98000_4000_M2 98000_6000_M2 0.022
r 98000_6000_M2 98000_8000_M2 0.022
r 98000_8000_M2 98000_10000_M2 0.022
r 98000_10000_M2 98000_12000_M2 0.022
r 98000_12000_M2 98000_14000_M2 0.022
r 98000_14000_M2 98000_16000_M2 0.022
r 98000_16000_M2 98000_18000_M2 0.022
r 98000_18000_M2 98000_20000_M2 0.022
r 98000_20000_M2 98000_22000_M2 0.022
r 98000_22000_M2 98000_24000_M2 0.022
r 98000_24000_M2 98000_26000_M2 0.022
r 98000_26000_M2 98000_28000_M2 0.022
r 98000_28000_M2 98000_30000_M2 0.022
r 98000_30000_M2 98000_32000_M2 0.022
r 98000_32000_M2 98000_34000_M2 0.022
r 98000_34000_M2 98000_36000_M2 0.022
r 98000_36000_M2 98000_38000_M2 0.022
r 98000_38000_M2 98000_40000_M2 0.022
r 98000_40000_M2 98000_42000_M2 0.022
r 98000_42000_M2 98000_44000_M2 0.022
r 98000_44000_M2 98000_46000_M2 0.022
r 98000_46000_M2 98000_48000_M2 0.022
r 98000_48000_M2 98000_50000_M2 0.022
r 98000_50000_M2 98000_52000_M2 0.022
r 98000_52000_M2 98000_54000_M2 0.022
r 98000_54000_M2 98000_56000_M2 0.022
r 98000_56000_M2 98000_58000_M2 0.022
r 98000_58000_M2 98000_60000_M2 0.022
r 98000_60000_M2 98000_62000_M2 0.022
r 98000_62000_M2 98000_64000_M2 0.022
r 98000_64000_M2 98000_66000_M2 0.022
r 98000_66000_M2 98000_68000_M2 0.022
r 98000_68000_M2 98000_70000_M2 0.022
r 98000_70000_M2 98000_72000_M2 0.022
r 98000_72000_M2 98000_74000_M2 0.022
r 98000_74000_M2 98000_76000_M2 0.022
r 98000_76000_M2 98000_78000_M2 0.022
r 98000_78000_M2 98000_80000_M2 0.022
r 98000_80000_M2 98000_82000_M2 0.022
r 98000_82000_M2 98000_84000_M2 0.022
r 98000_84000_M2 98000_86000_M2 0.022
r 98000_86000_M2 98000_88000_M2 0.022
r 98000_88000_M2 98000_90000_M2 0.022
r 98000_90000_M2 98000_92000_M2 0.022
r 98000_92000_M2 98000_94000_M2 0.022
r 98000_94000_M2 98000_96000_M2 0.022
r 98000_96000_M2 98000_98000_M2 0.022
r 98000_98000_M2 98000_100000_M2 0.022
r 100000_2000_M2 100000_4000_M2 0.022
r 100000_4000_M2 100000_6000_M2 0.022
r 100000_6000_M2 100000_8000_M2 0.022
r 100000_8000_M2 100000_10000_M2 0.022
r 100000_10000_M2 100000_12000_M2 0.022
r 100000_12000_M2 100000_14000_M2 0.022
r 100000_14000_M2 100000_16000_M2 0.022
r 100000_16000_M2 100000_18000_M2 0.022
r 100000_18000_M2 100000_20000_M2 0.022
r 100000_20000_M2 100000_22000_M2 0.022
r 100000_22000_M2 100000_24000_M2 0.022
r 100000_24000_M2 100000_26000_M2 0.022
r 100000_26000_M2 100000_28000_M2 0.022
r 100000_28000_M2 100000_30000_M2 0.022
r 100000_30000_M2 100000_32000_M2 0.022
r 100000_32000_M2 100000_34000_M2 0.022
r 100000_34000_M2 100000_36000_M2 0.022
r 100000_36000_M2 100000_38000_M2 0.022
r 100000_38000_M2 100000_40000_M2 0.022
r 100000_40000_M2 100000_42000_M2 0.022
r 100000_42000_M2 100000_44000_M2 0.022
r 100000_44000_M2 100000_46000_M2 0.022
r 100000_46000_M2 100000_48000_M2 0.022
r 100000_48000_M2 100000_50000_M2 0.022
r 100000_50000_M2 100000_52000_M2 0.022
r 100000_52000_M2 100000_54000_M2 0.022
r 100000_54000_M2 100000_56000_M2 0.022
r 100000_56000_M2 100000_58000_M2 0.022
r 100000_58000_M2 100000_60000_M2 0.022
r 100000_60000_M2 100000_62000_M2 0.022
r 100000_62000_M2 100000_64000_M2 0.022
r 100000_64000_M2 100000_66000_M2 0.022
r 100000_66000_M2 100000_68000_M2 0.022
r 100000_68000_M2 100000_70000_M2 0.022
r 100000_70000_M2 100000_72000_M2 0.022
r 100000_72000_M2 100000_74000_M2 0.022
r 100000_74000_M2 100000_76000_M2 0.022
r 100000_76000_M2 100000_78000_M2 0.022
r 100000_78000_M2 100000_80000_M2 0.022
r 100000_80000_M2 100000_82000_M2 0.022
r 100000_82000_M2 100000_84000_M2 0.022
r 100000_84000_M2 100000_86000_M2 0.022
r 100000_86000_M2 100000_88000_M2 0.022
r 100000_88000_M2 100000_90000_M2 0.022
r 100000_90000_M2 100000_92000_M2 0.022
r 100000_92000_M2 100000_94000_M2 0.022
r 100000_94000_M2 100000_96000_M2 0.022
r 100000_96000_M2 100000_98000_M2 0.022
r 100000_98000_M2 100000_100000_M2 0.022

* ============================================================================
* Layer M3 - 25x25 grid
* ============================================================================

* M3 Horizontal resistors
r 4000_4000_M3 8000_4000_M3 0.015
r 8000_4000_M3 12000_4000_M3 0.015
r 12000_4000_M3 16000_4000_M3 0.015
r 16000_4000_M3 20000_4000_M3 0.015
r 20000_4000_M3 24000_4000_M3 0.015
r 24000_4000_M3 28000_4000_M3 0.015
r 28000_4000_M3 32000_4000_M3 0.015
r 32000_4000_M3 36000_4000_M3 0.015
r 36000_4000_M3 40000_4000_M3 0.015
r 40000_4000_M3 44000_4000_M3 0.015
r 44000_4000_M3 48000_4000_M3 0.015
r 48000_4000_M3 52000_4000_M3 0.015
r 52000_4000_M3 56000_4000_M3 0.015
r 56000_4000_M3 60000_4000_M3 0.015
r 60000_4000_M3 64000_4000_M3 0.015
r 64000_4000_M3 68000_4000_M3 0.015
r 68000_4000_M3 72000_4000_M3 0.015
r 72000_4000_M3 76000_4000_M3 0.015
r 76000_4000_M3 80000_4000_M3 0.015
r 80000_4000_M3 84000_4000_M3 0.015
r 84000_4000_M3 88000_4000_M3 0.015
r 88000_4000_M3 92000_4000_M3 0.015
r 92000_4000_M3 96000_4000_M3 0.015
r 96000_4000_M3 100000_4000_M3 0.015
r 4000_8000_M3 8000_8000_M3 0.015
r 8000_8000_M3 12000_8000_M3 0.015
r 12000_8000_M3 16000_8000_M3 0.015
r 16000_8000_M3 20000_8000_M3 0.015
r 20000_8000_M3 24000_8000_M3 0.015
r 24000_8000_M3 28000_8000_M3 0.015
r 28000_8000_M3 32000_8000_M3 0.015
r 32000_8000_M3 36000_8000_M3 0.015
r 36000_8000_M3 40000_8000_M3 0.015
r 40000_8000_M3 44000_8000_M3 0.015
r 44000_8000_M3 48000_8000_M3 0.015
r 48000_8000_M3 52000_8000_M3 0.015
r 52000_8000_M3 56000_8000_M3 0.015
r 56000_8000_M3 60000_8000_M3 0.015
r 60000_8000_M3 64000_8000_M3 0.015
r 64000_8000_M3 68000_8000_M3 0.015
r 68000_8000_M3 72000_8000_M3 0.015
r 72000_8000_M3 76000_8000_M3 0.015
r 76000_8000_M3 80000_8000_M3 0.015
r 80000_8000_M3 84000_8000_M3 0.015
r 84000_8000_M3 88000_8000_M3 0.015
r 88000_8000_M3 92000_8000_M3 0.015
r 92000_8000_M3 96000_8000_M3 0.015
r 96000_8000_M3 100000_8000_M3 0.015
r 4000_12000_M3 8000_12000_M3 0.015
r 8000_12000_M3 12000_12000_M3 0.015
r 12000_12000_M3 16000_12000_M3 0.015
r 16000_12000_M3 20000_12000_M3 0.015
r 20000_12000_M3 24000_12000_M3 0.015
r 24000_12000_M3 28000_12000_M3 0.015
r 28000_12000_M3 32000_12000_M3 0.015
r 32000_12000_M3 36000_12000_M3 0.015
r 36000_12000_M3 40000_12000_M3 0.015
r 40000_12000_M3 44000_12000_M3 0.015
r 44000_12000_M3 48000_12000_M3 0.015
r 48000_12000_M3 52000_12000_M3 0.015
r 52000_12000_M3 56000_12000_M3 0.015
r 56000_12000_M3 60000_12000_M3 0.015
r 60000_12000_M3 64000_12000_M3 0.015
r 64000_12000_M3 68000_12000_M3 0.015
r 68000_12000_M3 72000_12000_M3 0.015
r 72000_12000_M3 76000_12000_M3 0.015
r 76000_12000_M3 80000_12000_M3 0.015
r 80000_12000_M3 84000_12000_M3 0.015
r 84000_12000_M3 88000_12000_M3 0.015
r 88000_12000_M3 92000_12000_M3 0.015
r 92000_12000_M3 96000_12000_M3 0.015
r 96000_12000_M3 100000_12000_M3 0.015
r 4000_16000_M3 8000_16000_M3 0.015
r 8000_16000_M3 12000_16000_M3 0.015
r 12000_16000_M3 16000_16000_M3 0.015
r 16000_16000_M3 20000_16000_M3 0.015
r 20000_16000_M3 24000_16000_M3 0.015
r 24000_16000_M3 28000_16000_M3 0.015
r 28000_16000_M3 32000_16000_M3 0.015
r 32000_16000_M3 36000_16000_M3 0.015
r 36000_16000_M3 40000_16000_M3 0.015
r 40000_16000_M3 44000_16000_M3 0.015
r 44000_16000_M3 48000_16000_M3 0.015
r 48000_16000_M3 52000_16000_M3 0.015
r 52000_16000_M3 56000_16000_M3 0.015
r 56000_16000_M3 60000_16000_M3 0.015
r 60000_16000_M3 64000_16000_M3 0.015
r 64000_16000_M3 68000_16000_M3 0.015
r 68000_16000_M3 72000_16000_M3 0.015
r 72000_16000_M3 76000_16000_M3 0.015
r 76000_16000_M3 80000_16000_M3 0.015
r 80000_16000_M3 84000_16000_M3 0.015
r 84000_16000_M3 88000_16000_M3 0.015
r 88000_16000_M3 92000_16000_M3 0.015
r 92000_16000_M3 96000_16000_M3 0.015
r 96000_16000_M3 100000_16000_M3 0.015
r 4000_20000_M3 8000_20000_M3 0.015
r 8000_20000_M3 12000_20000_M3 0.015
r 12000_20000_M3 16000_20000_M3 0.015
r 16000_20000_M3 20000_20000_M3 0.015
r 20000_20000_M3 24000_20000_M3 0.015
r 24000_20000_M3 28000_20000_M3 0.015
r 28000_20000_M3 32000_20000_M3 0.015
r 32000_20000_M3 36000_20000_M3 0.015
r 36000_20000_M3 40000_20000_M3 0.015
r 40000_20000_M3 44000_20000_M3 0.015
r 44000_20000_M3 48000_20000_M3 0.015
r 48000_20000_M3 52000_20000_M3 0.015
r 52000_20000_M3 56000_20000_M3 0.015
r 56000_20000_M3 60000_20000_M3 0.015
r 60000_20000_M3 64000_20000_M3 0.015
r 64000_20000_M3 68000_20000_M3 0.015
r 68000_20000_M3 72000_20000_M3 0.015
r 72000_20000_M3 76000_20000_M3 0.015
r 76000_20000_M3 80000_20000_M3 0.015
r 80000_20000_M3 84000_20000_M3 0.015
r 84000_20000_M3 88000_20000_M3 0.015
r 88000_20000_M3 92000_20000_M3 0.015
r 92000_20000_M3 96000_20000_M3 0.015
r 96000_20000_M3 100000_20000_M3 0.015
r 4000_24000_M3 8000_24000_M3 0.015
r 8000_24000_M3 12000_24000_M3 0.015
r 12000_24000_M3 16000_24000_M3 0.015
r 16000_24000_M3 20000_24000_M3 0.015
r 20000_24000_M3 24000_24000_M3 0.015
r 24000_24000_M3 28000_24000_M3 0.015
r 28000_24000_M3 32000_24000_M3 0.015
r 32000_24000_M3 36000_24000_M3 0.015
r 36000_24000_M3 40000_24000_M3 0.015
r 40000_24000_M3 44000_24000_M3 0.015
r 44000_24000_M3 48000_24000_M3 0.015
r 48000_24000_M3 52000_24000_M3 0.015
r 52000_24000_M3 56000_24000_M3 0.015
r 56000_24000_M3 60000_24000_M3 0.015
r 60000_24000_M3 64000_24000_M3 0.015
r 64000_24000_M3 68000_24000_M3 0.015
r 68000_24000_M3 72000_24000_M3 0.015
r 72000_24000_M3 76000_24000_M3 0.015
r 76000_24000_M3 80000_24000_M3 0.015
r 80000_24000_M3 84000_24000_M3 0.015
r 84000_24000_M3 88000_24000_M3 0.015
r 88000_24000_M3 92000_24000_M3 0.015
r 92000_24000_M3 96000_24000_M3 0.015
r 96000_24000_M3 100000_24000_M3 0.015
r 4000_28000_M3 8000_28000_M3 0.015
r 8000_28000_M3 12000_28000_M3 0.015
r 12000_28000_M3 16000_28000_M3 0.015
r 16000_28000_M3 20000_28000_M3 0.015
r 20000_28000_M3 24000_28000_M3 0.015
r 24000_28000_M3 28000_28000_M3 0.015
r 28000_28000_M3 32000_28000_M3 0.015
r 32000_28000_M3 36000_28000_M3 0.015
r 36000_28000_M3 40000_28000_M3 0.015
r 40000_28000_M3 44000_28000_M3 0.015
r 44000_28000_M3 48000_28000_M3 0.015
r 48000_28000_M3 52000_28000_M3 0.015
r 52000_28000_M3 56000_28000_M3 0.015
r 56000_28000_M3 60000_28000_M3 0.015
r 60000_28000_M3 64000_28000_M3 0.015
r 64000_28000_M3 68000_28000_M3 0.015
r 68000_28000_M3 72000_28000_M3 0.015
r 72000_28000_M3 76000_28000_M3 0.015
r 76000_28000_M3 80000_28000_M3 0.015
r 80000_28000_M3 84000_28000_M3 0.015
r 84000_28000_M3 88000_28000_M3 0.015
r 88000_28000_M3 92000_28000_M3 0.015
r 92000_28000_M3 96000_28000_M3 0.015
r 96000_28000_M3 100000_28000_M3 0.015
r 4000_32000_M3 8000_32000_M3 0.015
r 8000_32000_M3 12000_32000_M3 0.015
r 12000_32000_M3 16000_32000_M3 0.015
r 16000_32000_M3 20000_32000_M3 0.015
r 20000_32000_M3 24000_32000_M3 0.015
r 24000_32000_M3 28000_32000_M3 0.015
r 28000_32000_M3 32000_32000_M3 0.015
r 32000_32000_M3 36000_32000_M3 0.015
r 36000_32000_M3 40000_32000_M3 0.015
r 40000_32000_M3 44000_32000_M3 0.015
r 44000_32000_M3 48000_32000_M3 0.015
r 48000_32000_M3 52000_32000_M3 0.015
r 52000_32000_M3 56000_32000_M3 0.015
r 56000_32000_M3 60000_32000_M3 0.015
r 60000_32000_M3 64000_32000_M3 0.015
r 64000_32000_M3 68000_32000_M3 0.015
r 68000_32000_M3 72000_32000_M3 0.015
r 72000_32000_M3 76000_32000_M3 0.015
r 76000_32000_M3 80000_32000_M3 0.015
r 80000_32000_M3 84000_32000_M3 0.015
r 84000_32000_M3 88000_32000_M3 0.015
r 88000_32000_M3 92000_32000_M3 0.015
r 92000_32000_M3 96000_32000_M3 0.015
r 96000_32000_M3 100000_32000_M3 0.015
r 4000_36000_M3 8000_36000_M3 0.015
r 8000_36000_M3 12000_36000_M3 0.015
r 12000_36000_M3 16000_36000_M3 0.015
r 16000_36000_M3 20000_36000_M3 0.015
r 20000_36000_M3 24000_36000_M3 0.015
r 24000_36000_M3 28000_36000_M3 0.015
r 28000_36000_M3 32000_36000_M3 0.015
r 32000_36000_M3 36000_36000_M3 0.015
r 36000_36000_M3 40000_36000_M3 0.015
r 40000_36000_M3 44000_36000_M3 0.015
r 44000_36000_M3 48000_36000_M3 0.015
r 48000_36000_M3 52000_36000_M3 0.015
r 52000_36000_M3 56000_36000_M3 0.015
r 56000_36000_M3 60000_36000_M3 0.015
r 60000_36000_M3 64000_36000_M3 0.015
r 64000_36000_M3 68000_36000_M3 0.015
r 68000_36000_M3 72000_36000_M3 0.015
r 72000_36000_M3 76000_36000_M3 0.015
r 76000_36000_M3 80000_36000_M3 0.015
r 80000_36000_M3 84000_36000_M3 0.015
r 84000_36000_M3 88000_36000_M3 0.015
r 88000_36000_M3 92000_36000_M3 0.015
r 92000_36000_M3 96000_36000_M3 0.015
r 96000_36000_M3 100000_36000_M3 0.015
r 4000_40000_M3 8000_40000_M3 0.015
r 8000_40000_M3 12000_40000_M3 0.015
r 12000_40000_M3 16000_40000_M3 0.015
r 16000_40000_M3 20000_40000_M3 0.015
r 20000_40000_M3 24000_40000_M3 0.015
r 24000_40000_M3 28000_40000_M3 0.015
r 28000_40000_M3 32000_40000_M3 0.015
r 32000_40000_M3 36000_40000_M3 0.015
r 36000_40000_M3 40000_40000_M3 0.015
r 40000_40000_M3 44000_40000_M3 0.015
r 44000_40000_M3 48000_40000_M3 0.015
r 48000_40000_M3 52000_40000_M3 0.015
r 52000_40000_M3 56000_40000_M3 0.015
r 56000_40000_M3 60000_40000_M3 0.015
r 60000_40000_M3 64000_40000_M3 0.015
r 64000_40000_M3 68000_40000_M3 0.015
r 68000_40000_M3 72000_40000_M3 0.015
r 72000_40000_M3 76000_40000_M3 0.015
r 76000_40000_M3 80000_40000_M3 0.015
r 80000_40000_M3 84000_40000_M3 0.015
r 84000_40000_M3 88000_40000_M3 0.015
r 88000_40000_M3 92000_40000_M3 0.015
r 92000_40000_M3 96000_40000_M3 0.015
r 96000_40000_M3 100000_40000_M3 0.015
r 4000_44000_M3 8000_44000_M3 0.015
r 8000_44000_M3 12000_44000_M3 0.015
r 12000_44000_M3 16000_44000_M3 0.015
r 16000_44000_M3 20000_44000_M3 0.015
r 20000_44000_M3 24000_44000_M3 0.015
r 24000_44000_M3 28000_44000_M3 0.015
r 28000_44000_M3 32000_44000_M3 0.015
r 32000_44000_M3 36000_44000_M3 0.015
r 36000_44000_M3 40000_44000_M3 0.015
r 40000_44000_M3 44000_44000_M3 0.015
r 44000_44000_M3 48000_44000_M3 0.015
r 48000_44000_M3 52000_44000_M3 0.015
r 52000_44000_M3 56000_44000_M3 0.015
r 56000_44000_M3 60000_44000_M3 0.015
r 60000_44000_M3 64000_44000_M3 0.015
r 64000_44000_M3 68000_44000_M3 0.015
r 68000_44000_M3 72000_44000_M3 0.015
r 72000_44000_M3 76000_44000_M3 0.015
r 76000_44000_M3 80000_44000_M3 0.015
r 80000_44000_M3 84000_44000_M3 0.015
r 84000_44000_M3 88000_44000_M3 0.015
r 88000_44000_M3 92000_44000_M3 0.015
r 92000_44000_M3 96000_44000_M3 0.015
r 96000_44000_M3 100000_44000_M3 0.015
r 4000_48000_M3 8000_48000_M3 0.015
r 8000_48000_M3 12000_48000_M3 0.015
r 12000_48000_M3 16000_48000_M3 0.015
r 16000_48000_M3 20000_48000_M3 0.015
r 20000_48000_M3 24000_48000_M3 0.015
r 24000_48000_M3 28000_48000_M3 0.015
r 28000_48000_M3 32000_48000_M3 0.015
r 32000_48000_M3 36000_48000_M3 0.015
r 36000_48000_M3 40000_48000_M3 0.015
r 40000_48000_M3 44000_48000_M3 0.015
r 44000_48000_M3 48000_48000_M3 0.015
r 48000_48000_M3 52000_48000_M3 0.015
r 52000_48000_M3 56000_48000_M3 0.015
r 56000_48000_M3 60000_48000_M3 0.015
r 60000_48000_M3 64000_48000_M3 0.015
r 64000_48000_M3 68000_48000_M3 0.015
r 68000_48000_M3 72000_48000_M3 0.015
r 72000_48000_M3 76000_48000_M3 0.015
r 76000_48000_M3 80000_48000_M3 0.015
r 80000_48000_M3 84000_48000_M3 0.015
r 84000_48000_M3 88000_48000_M3 0.015
r 88000_48000_M3 92000_48000_M3 0.015
r 92000_48000_M3 96000_48000_M3 0.015
r 96000_48000_M3 100000_48000_M3 0.015
r 4000_52000_M3 8000_52000_M3 0.015
r 8000_52000_M3 12000_52000_M3 0.015
r 12000_52000_M3 16000_52000_M3 0.015
r 16000_52000_M3 20000_52000_M3 0.015
r 20000_52000_M3 24000_52000_M3 0.015
r 24000_52000_M3 28000_52000_M3 0.015
r 28000_52000_M3 32000_52000_M3 0.015
r 32000_52000_M3 36000_52000_M3 0.015
r 36000_52000_M3 40000_52000_M3 0.015
r 40000_52000_M3 44000_52000_M3 0.015
r 44000_52000_M3 48000_52000_M3 0.015
r 48000_52000_M3 52000_52000_M3 0.015
r 52000_52000_M3 56000_52000_M3 0.015
r 56000_52000_M3 60000_52000_M3 0.015
r 60000_52000_M3 64000_52000_M3 0.015
r 64000_52000_M3 68000_52000_M3 0.015
r 68000_52000_M3 72000_52000_M3 0.015
r 72000_52000_M3 76000_52000_M3 0.015
r 76000_52000_M3 80000_52000_M3 0.015
r 80000_52000_M3 84000_52000_M3 0.015
r 84000_52000_M3 88000_52000_M3 0.015
r 88000_52000_M3 92000_52000_M3 0.015
r 92000_52000_M3 96000_52000_M3 0.015
r 96000_52000_M3 100000_52000_M3 0.015
r 4000_56000_M3 8000_56000_M3 0.015
r 8000_56000_M3 12000_56000_M3 0.015
r 12000_56000_M3 16000_56000_M3 0.015
r 16000_56000_M3 20000_56000_M3 0.015
r 20000_56000_M3 24000_56000_M3 0.015
r 24000_56000_M3 28000_56000_M3 0.015
r 28000_56000_M3 32000_56000_M3 0.015
r 32000_56000_M3 36000_56000_M3 0.015
r 36000_56000_M3 40000_56000_M3 0.015
r 40000_56000_M3 44000_56000_M3 0.015
r 44000_56000_M3 48000_56000_M3 0.015
r 48000_56000_M3 52000_56000_M3 0.015
r 52000_56000_M3 56000_56000_M3 0.015
r 56000_56000_M3 60000_56000_M3 0.015
r 60000_56000_M3 64000_56000_M3 0.015
r 64000_56000_M3 68000_56000_M3 0.015
r 68000_56000_M3 72000_56000_M3 0.015
r 72000_56000_M3 76000_56000_M3 0.015
r 76000_56000_M3 80000_56000_M3 0.015
r 80000_56000_M3 84000_56000_M3 0.015
r 84000_56000_M3 88000_56000_M3 0.015
r 88000_56000_M3 92000_56000_M3 0.015
r 92000_56000_M3 96000_56000_M3 0.015
r 96000_56000_M3 100000_56000_M3 0.015
r 4000_60000_M3 8000_60000_M3 0.015
r 8000_60000_M3 12000_60000_M3 0.015
r 12000_60000_M3 16000_60000_M3 0.015
r 16000_60000_M3 20000_60000_M3 0.015
r 20000_60000_M3 24000_60000_M3 0.015
r 24000_60000_M3 28000_60000_M3 0.015
r 28000_60000_M3 32000_60000_M3 0.015
r 32000_60000_M3 36000_60000_M3 0.015
r 36000_60000_M3 40000_60000_M3 0.015
r 40000_60000_M3 44000_60000_M3 0.015
r 44000_60000_M3 48000_60000_M3 0.015
r 48000_60000_M3 52000_60000_M3 0.015
r 52000_60000_M3 56000_60000_M3 0.015
r 56000_60000_M3 60000_60000_M3 0.015
r 60000_60000_M3 64000_60000_M3 0.015
r 64000_60000_M3 68000_60000_M3 0.015
r 68000_60000_M3 72000_60000_M3 0.015
r 72000_60000_M3 76000_60000_M3 0.015
r 76000_60000_M3 80000_60000_M3 0.015
r 80000_60000_M3 84000_60000_M3 0.015
r 84000_60000_M3 88000_60000_M3 0.015
r 88000_60000_M3 92000_60000_M3 0.015
r 92000_60000_M3 96000_60000_M3 0.015
r 96000_60000_M3 100000_60000_M3 0.015
r 4000_64000_M3 8000_64000_M3 0.015
r 8000_64000_M3 12000_64000_M3 0.015
r 12000_64000_M3 16000_64000_M3 0.015
r 16000_64000_M3 20000_64000_M3 0.015
r 20000_64000_M3 24000_64000_M3 0.015
r 24000_64000_M3 28000_64000_M3 0.015
r 28000_64000_M3 32000_64000_M3 0.015
r 32000_64000_M3 36000_64000_M3 0.015
r 36000_64000_M3 40000_64000_M3 0.015
r 40000_64000_M3 44000_64000_M3 0.015
r 44000_64000_M3 48000_64000_M3 0.015
r 48000_64000_M3 52000_64000_M3 0.015
r 52000_64000_M3 56000_64000_M3 0.015
r 56000_64000_M3 60000_64000_M3 0.015
r 60000_64000_M3 64000_64000_M3 0.015
r 64000_64000_M3 68000_64000_M3 0.015
r 68000_64000_M3 72000_64000_M3 0.015
r 72000_64000_M3 76000_64000_M3 0.015
r 76000_64000_M3 80000_64000_M3 0.015
r 80000_64000_M3 84000_64000_M3 0.015
r 84000_64000_M3 88000_64000_M3 0.015
r 88000_64000_M3 92000_64000_M3 0.015
r 92000_64000_M3 96000_64000_M3 0.015
r 96000_64000_M3 100000_64000_M3 0.015
r 4000_68000_M3 8000_68000_M3 0.015
r 8000_68000_M3 12000_68000_M3 0.015
r 12000_68000_M3 16000_68000_M3 0.015
r 16000_68000_M3 20000_68000_M3 0.015
r 20000_68000_M3 24000_68000_M3 0.015
r 24000_68000_M3 28000_68000_M3 0.015
r 28000_68000_M3 32000_68000_M3 0.015
r 32000_68000_M3 36000_68000_M3 0.015
r 36000_68000_M3 40000_68000_M3 0.015
r 40000_68000_M3 44000_68000_M3 0.015
r 44000_68000_M3 48000_68000_M3 0.015
r 48000_68000_M3 52000_68000_M3 0.015
r 52000_68000_M3 56000_68000_M3 0.015
r 56000_68000_M3 60000_68000_M3 0.015
r 60000_68000_M3 64000_68000_M3 0.015
r 64000_68000_M3 68000_68000_M3 0.015
r 68000_68000_M3 72000_68000_M3 0.015
r 72000_68000_M3 76000_68000_M3 0.015
r 76000_68000_M3 80000_68000_M3 0.015
r 80000_68000_M3 84000_68000_M3 0.015
r 84000_68000_M3 88000_68000_M3 0.015
r 88000_68000_M3 92000_68000_M3 0.015
r 92000_68000_M3 96000_68000_M3 0.015
r 96000_68000_M3 100000_68000_M3 0.015
r 4000_72000_M3 8000_72000_M3 0.015
r 8000_72000_M3 12000_72000_M3 0.015
r 12000_72000_M3 16000_72000_M3 0.015
r 16000_72000_M3 20000_72000_M3 0.015
r 20000_72000_M3 24000_72000_M3 0.015
r 24000_72000_M3 28000_72000_M3 0.015
r 28000_72000_M3 32000_72000_M3 0.015
r 32000_72000_M3 36000_72000_M3 0.015
r 36000_72000_M3 40000_72000_M3 0.015
r 40000_72000_M3 44000_72000_M3 0.015
r 44000_72000_M3 48000_72000_M3 0.015
r 48000_72000_M3 52000_72000_M3 0.015
r 52000_72000_M3 56000_72000_M3 0.015
r 56000_72000_M3 60000_72000_M3 0.015
r 60000_72000_M3 64000_72000_M3 0.015
r 64000_72000_M3 68000_72000_M3 0.015
r 68000_72000_M3 72000_72000_M3 0.015
r 72000_72000_M3 76000_72000_M3 0.015
r 76000_72000_M3 80000_72000_M3 0.015
r 80000_72000_M3 84000_72000_M3 0.015
r 84000_72000_M3 88000_72000_M3 0.015
r 88000_72000_M3 92000_72000_M3 0.015
r 92000_72000_M3 96000_72000_M3 0.015
r 96000_72000_M3 100000_72000_M3 0.015
r 4000_76000_M3 8000_76000_M3 0.015
r 8000_76000_M3 12000_76000_M3 0.015
r 12000_76000_M3 16000_76000_M3 0.015
r 16000_76000_M3 20000_76000_M3 0.015
r 20000_76000_M3 24000_76000_M3 0.015
r 24000_76000_M3 28000_76000_M3 0.015
r 28000_76000_M3 32000_76000_M3 0.015
r 32000_76000_M3 36000_76000_M3 0.015
r 36000_76000_M3 40000_76000_M3 0.015
r 40000_76000_M3 44000_76000_M3 0.015
r 44000_76000_M3 48000_76000_M3 0.015
r 48000_76000_M3 52000_76000_M3 0.015
r 52000_76000_M3 56000_76000_M3 0.015
r 56000_76000_M3 60000_76000_M3 0.015
r 60000_76000_M3 64000_76000_M3 0.015
r 64000_76000_M3 68000_76000_M3 0.015
r 68000_76000_M3 72000_76000_M3 0.015
r 72000_76000_M3 76000_76000_M3 0.015
r 76000_76000_M3 80000_76000_M3 0.015
r 80000_76000_M3 84000_76000_M3 0.015
r 84000_76000_M3 88000_76000_M3 0.015
r 88000_76000_M3 92000_76000_M3 0.015
r 92000_76000_M3 96000_76000_M3 0.015
r 96000_76000_M3 100000_76000_M3 0.015
r 4000_80000_M3 8000_80000_M3 0.015
r 8000_80000_M3 12000_80000_M3 0.015
r 12000_80000_M3 16000_80000_M3 0.015
r 16000_80000_M3 20000_80000_M3 0.015
r 20000_80000_M3 24000_80000_M3 0.015
r 24000_80000_M3 28000_80000_M3 0.015
r 28000_80000_M3 32000_80000_M3 0.015
r 32000_80000_M3 36000_80000_M3 0.015
r 36000_80000_M3 40000_80000_M3 0.015
r 40000_80000_M3 44000_80000_M3 0.015
r 44000_80000_M3 48000_80000_M3 0.015
r 48000_80000_M3 52000_80000_M3 0.015
r 52000_80000_M3 56000_80000_M3 0.015
r 56000_80000_M3 60000_80000_M3 0.015
r 60000_80000_M3 64000_80000_M3 0.015
r 64000_80000_M3 68000_80000_M3 0.015
r 68000_80000_M3 72000_80000_M3 0.015
r 72000_80000_M3 76000_80000_M3 0.015
r 76000_80000_M3 80000_80000_M3 0.015
r 80000_80000_M3 84000_80000_M3 0.015
r 84000_80000_M3 88000_80000_M3 0.015
r 88000_80000_M3 92000_80000_M3 0.015
r 92000_80000_M3 96000_80000_M3 0.015
r 96000_80000_M3 100000_80000_M3 0.015
r 4000_84000_M3 8000_84000_M3 0.015
r 8000_84000_M3 12000_84000_M3 0.015
r 12000_84000_M3 16000_84000_M3 0.015
r 16000_84000_M3 20000_84000_M3 0.015
r 20000_84000_M3 24000_84000_M3 0.015
r 24000_84000_M3 28000_84000_M3 0.015
r 28000_84000_M3 32000_84000_M3 0.015
r 32000_84000_M3 36000_84000_M3 0.015
r 36000_84000_M3 40000_84000_M3 0.015
r 40000_84000_M3 44000_84000_M3 0.015
r 44000_84000_M3 48000_84000_M3 0.015
r 48000_84000_M3 52000_84000_M3 0.015
r 52000_84000_M3 56000_84000_M3 0.015
r 56000_84000_M3 60000_84000_M3 0.015
r 60000_84000_M3 64000_84000_M3 0.015
r 64000_84000_M3 68000_84000_M3 0.015
r 68000_84000_M3 72000_84000_M3 0.015
r 72000_84000_M3 76000_84000_M3 0.015
r 76000_84000_M3 80000_84000_M3 0.015
r 80000_84000_M3 84000_84000_M3 0.015
r 84000_84000_M3 88000_84000_M3 0.015
r 88000_84000_M3 92000_84000_M3 0.015
r 92000_84000_M3 96000_84000_M3 0.015
r 96000_84000_M3 100000_84000_M3 0.015
r 4000_88000_M3 8000_88000_M3 0.015
r 8000_88000_M3 12000_88000_M3 0.015
r 12000_88000_M3 16000_88000_M3 0.015
r 16000_88000_M3 20000_88000_M3 0.015
r 20000_88000_M3 24000_88000_M3 0.015
r 24000_88000_M3 28000_88000_M3 0.015
r 28000_88000_M3 32000_88000_M3 0.015
r 32000_88000_M3 36000_88000_M3 0.015
r 36000_88000_M3 40000_88000_M3 0.015
r 40000_88000_M3 44000_88000_M3 0.015
r 44000_88000_M3 48000_88000_M3 0.015
r 48000_88000_M3 52000_88000_M3 0.015
r 52000_88000_M3 56000_88000_M3 0.015
r 56000_88000_M3 60000_88000_M3 0.015
r 60000_88000_M3 64000_88000_M3 0.015
r 64000_88000_M3 68000_88000_M3 0.015
r 68000_88000_M3 72000_88000_M3 0.015
r 72000_88000_M3 76000_88000_M3 0.015
r 76000_88000_M3 80000_88000_M3 0.015
r 80000_88000_M3 84000_88000_M3 0.015
r 84000_88000_M3 88000_88000_M3 0.015
r 88000_88000_M3 92000_88000_M3 0.015
r 92000_88000_M3 96000_88000_M3 0.015
r 96000_88000_M3 100000_88000_M3 0.015
r 4000_92000_M3 8000_92000_M3 0.015
r 8000_92000_M3 12000_92000_M3 0.015
r 12000_92000_M3 16000_92000_M3 0.015
r 16000_92000_M3 20000_92000_M3 0.015
r 20000_92000_M3 24000_92000_M3 0.015
r 24000_92000_M3 28000_92000_M3 0.015
r 28000_92000_M3 32000_92000_M3 0.015
r 32000_92000_M3 36000_92000_M3 0.015
r 36000_92000_M3 40000_92000_M3 0.015
r 40000_92000_M3 44000_92000_M3 0.015
r 44000_92000_M3 48000_92000_M3 0.015
r 48000_92000_M3 52000_92000_M3 0.015
r 52000_92000_M3 56000_92000_M3 0.015
r 56000_92000_M3 60000_92000_M3 0.015
r 60000_92000_M3 64000_92000_M3 0.015
r 64000_92000_M3 68000_92000_M3 0.015
r 68000_92000_M3 72000_92000_M3 0.015
r 72000_92000_M3 76000_92000_M3 0.015
r 76000_92000_M3 80000_92000_M3 0.015
r 80000_92000_M3 84000_92000_M3 0.015
r 84000_92000_M3 88000_92000_M3 0.015
r 88000_92000_M3 92000_92000_M3 0.015
r 92000_92000_M3 96000_92000_M3 0.015
r 96000_92000_M3 100000_92000_M3 0.015
r 4000_96000_M3 8000_96000_M3 0.015
r 8000_96000_M3 12000_96000_M3 0.015
r 12000_96000_M3 16000_96000_M3 0.015
r 16000_96000_M3 20000_96000_M3 0.015
r 20000_96000_M3 24000_96000_M3 0.015
r 24000_96000_M3 28000_96000_M3 0.015
r 28000_96000_M3 32000_96000_M3 0.015
r 32000_96000_M3 36000_96000_M3 0.015
r 36000_96000_M3 40000_96000_M3 0.015
r 40000_96000_M3 44000_96000_M3 0.015
r 44000_96000_M3 48000_96000_M3 0.015
r 48000_96000_M3 52000_96000_M3 0.015
r 52000_96000_M3 56000_96000_M3 0.015
r 56000_96000_M3 60000_96000_M3 0.015
r 60000_96000_M3 64000_96000_M3 0.015
r 64000_96000_M3 68000_96000_M3 0.015
r 68000_96000_M3 72000_96000_M3 0.015
r 72000_96000_M3 76000_96000_M3 0.015
r 76000_96000_M3 80000_96000_M3 0.015
r 80000_96000_M3 84000_96000_M3 0.015
r 84000_96000_M3 88000_96000_M3 0.015
r 88000_96000_M3 92000_96000_M3 0.015
r 92000_96000_M3 96000_96000_M3 0.015
r 96000_96000_M3 100000_96000_M3 0.015
r 4000_100000_M3 8000_100000_M3 0.015
r 8000_100000_M3 12000_100000_M3 0.015
r 12000_100000_M3 16000_100000_M3 0.015
r 16000_100000_M3 20000_100000_M3 0.015
r 20000_100000_M3 24000_100000_M3 0.015
r 24000_100000_M3 28000_100000_M3 0.015
r 28000_100000_M3 32000_100000_M3 0.015
r 32000_100000_M3 36000_100000_M3 0.015
r 36000_100000_M3 40000_100000_M3 0.015
r 40000_100000_M3 44000_100000_M3 0.015
r 44000_100000_M3 48000_100000_M3 0.015
r 48000_100000_M3 52000_100000_M3 0.015
r 52000_100000_M3 56000_100000_M3 0.015
r 56000_100000_M3 60000_100000_M3 0.015
r 60000_100000_M3 64000_100000_M3 0.015
r 64000_100000_M3 68000_100000_M3 0.015
r 68000_100000_M3 72000_100000_M3 0.015
r 72000_100000_M3 76000_100000_M3 0.015
r 76000_100000_M3 80000_100000_M3 0.015
r 80000_100000_M3 84000_100000_M3 0.015
r 84000_100000_M3 88000_100000_M3 0.015
r 88000_100000_M3 92000_100000_M3 0.015
r 92000_100000_M3 96000_100000_M3 0.015
r 96000_100000_M3 100000_100000_M3 0.015

* M3 Vertical resistors
r 4000_4000_M3 4000_8000_M3 0.018
r 4000_8000_M3 4000_12000_M3 0.018
r 4000_12000_M3 4000_16000_M3 0.018
r 4000_16000_M3 4000_20000_M3 0.018
r 4000_20000_M3 4000_24000_M3 0.018
r 4000_24000_M3 4000_28000_M3 0.018
r 4000_28000_M3 4000_32000_M3 0.018
r 4000_32000_M3 4000_36000_M3 0.018
r 4000_36000_M3 4000_40000_M3 0.018
r 4000_40000_M3 4000_44000_M3 0.018
r 4000_44000_M3 4000_48000_M3 0.018
r 4000_48000_M3 4000_52000_M3 0.018
r 4000_52000_M3 4000_56000_M3 0.018
r 4000_56000_M3 4000_60000_M3 0.018
r 4000_60000_M3 4000_64000_M3 0.018
r 4000_64000_M3 4000_68000_M3 0.018
r 4000_68000_M3 4000_72000_M3 0.018
r 4000_72000_M3 4000_76000_M3 0.018
r 4000_76000_M3 4000_80000_M3 0.018
r 4000_80000_M3 4000_84000_M3 0.018
r 4000_84000_M3 4000_88000_M3 0.018
r 4000_88000_M3 4000_92000_M3 0.018
r 4000_92000_M3 4000_96000_M3 0.018
r 4000_96000_M3 4000_100000_M3 0.018
r 8000_4000_M3 8000_8000_M3 0.018
r 8000_8000_M3 8000_12000_M3 0.018
r 8000_12000_M3 8000_16000_M3 0.018
r 8000_16000_M3 8000_20000_M3 0.018
r 8000_20000_M3 8000_24000_M3 0.018
r 8000_24000_M3 8000_28000_M3 0.018
r 8000_28000_M3 8000_32000_M3 0.018
r 8000_32000_M3 8000_36000_M3 0.018
r 8000_36000_M3 8000_40000_M3 0.018
r 8000_40000_M3 8000_44000_M3 0.018
r 8000_44000_M3 8000_48000_M3 0.018
r 8000_48000_M3 8000_52000_M3 0.018
r 8000_52000_M3 8000_56000_M3 0.018
r 8000_56000_M3 8000_60000_M3 0.018
r 8000_60000_M3 8000_64000_M3 0.018
r 8000_64000_M3 8000_68000_M3 0.018
r 8000_68000_M3 8000_72000_M3 0.018
r 8000_72000_M3 8000_76000_M3 0.018
r 8000_76000_M3 8000_80000_M3 0.018
r 8000_80000_M3 8000_84000_M3 0.018
r 8000_84000_M3 8000_88000_M3 0.018
r 8000_88000_M3 8000_92000_M3 0.018
r 8000_92000_M3 8000_96000_M3 0.018
r 8000_96000_M3 8000_100000_M3 0.018
r 12000_4000_M3 12000_8000_M3 0.018
r 12000_8000_M3 12000_12000_M3 0.018
r 12000_12000_M3 12000_16000_M3 0.018
r 12000_16000_M3 12000_20000_M3 0.018
r 12000_20000_M3 12000_24000_M3 0.018
r 12000_24000_M3 12000_28000_M3 0.018
r 12000_28000_M3 12000_32000_M3 0.018
r 12000_32000_M3 12000_36000_M3 0.018
r 12000_36000_M3 12000_40000_M3 0.018
r 12000_40000_M3 12000_44000_M3 0.018
r 12000_44000_M3 12000_48000_M3 0.018
r 12000_48000_M3 12000_52000_M3 0.018
r 12000_52000_M3 12000_56000_M3 0.018
r 12000_56000_M3 12000_60000_M3 0.018
r 12000_60000_M3 12000_64000_M3 0.018
r 12000_64000_M3 12000_68000_M3 0.018
r 12000_68000_M3 12000_72000_M3 0.018
r 12000_72000_M3 12000_76000_M3 0.018
r 12000_76000_M3 12000_80000_M3 0.018
r 12000_80000_M3 12000_84000_M3 0.018
r 12000_84000_M3 12000_88000_M3 0.018
r 12000_88000_M3 12000_92000_M3 0.018
r 12000_92000_M3 12000_96000_M3 0.018
r 12000_96000_M3 12000_100000_M3 0.018
r 16000_4000_M3 16000_8000_M3 0.018
r 16000_8000_M3 16000_12000_M3 0.018
r 16000_12000_M3 16000_16000_M3 0.018
r 16000_16000_M3 16000_20000_M3 0.018
r 16000_20000_M3 16000_24000_M3 0.018
r 16000_24000_M3 16000_28000_M3 0.018
r 16000_28000_M3 16000_32000_M3 0.018
r 16000_32000_M3 16000_36000_M3 0.018
r 16000_36000_M3 16000_40000_M3 0.018
r 16000_40000_M3 16000_44000_M3 0.018
r 16000_44000_M3 16000_48000_M3 0.018
r 16000_48000_M3 16000_52000_M3 0.018
r 16000_52000_M3 16000_56000_M3 0.018
r 16000_56000_M3 16000_60000_M3 0.018
r 16000_60000_M3 16000_64000_M3 0.018
r 16000_64000_M3 16000_68000_M3 0.018
r 16000_68000_M3 16000_72000_M3 0.018
r 16000_72000_M3 16000_76000_M3 0.018
r 16000_76000_M3 16000_80000_M3 0.018
r 16000_80000_M3 16000_84000_M3 0.018
r 16000_84000_M3 16000_88000_M3 0.018
r 16000_88000_M3 16000_92000_M3 0.018
r 16000_92000_M3 16000_96000_M3 0.018
r 16000_96000_M3 16000_100000_M3 0.018
r 20000_4000_M3 20000_8000_M3 0.018
r 20000_8000_M3 20000_12000_M3 0.018
r 20000_12000_M3 20000_16000_M3 0.018
r 20000_16000_M3 20000_20000_M3 0.018
r 20000_20000_M3 20000_24000_M3 0.018
r 20000_24000_M3 20000_28000_M3 0.018
r 20000_28000_M3 20000_32000_M3 0.018
r 20000_32000_M3 20000_36000_M3 0.018
r 20000_36000_M3 20000_40000_M3 0.018
r 20000_40000_M3 20000_44000_M3 0.018
r 20000_44000_M3 20000_48000_M3 0.018
r 20000_48000_M3 20000_52000_M3 0.018
r 20000_52000_M3 20000_56000_M3 0.018
r 20000_56000_M3 20000_60000_M3 0.018
r 20000_60000_M3 20000_64000_M3 0.018
r 20000_64000_M3 20000_68000_M3 0.018
r 20000_68000_M3 20000_72000_M3 0.018
r 20000_72000_M3 20000_76000_M3 0.018
r 20000_76000_M3 20000_80000_M3 0.018
r 20000_80000_M3 20000_84000_M3 0.018
r 20000_84000_M3 20000_88000_M3 0.018
r 20000_88000_M3 20000_92000_M3 0.018
r 20000_92000_M3 20000_96000_M3 0.018
r 20000_96000_M3 20000_100000_M3 0.018
r 24000_4000_M3 24000_8000_M3 0.018
r 24000_8000_M3 24000_12000_M3 0.018
r 24000_12000_M3 24000_16000_M3 0.018
r 24000_16000_M3 24000_20000_M3 0.018
r 24000_20000_M3 24000_24000_M3 0.018
r 24000_24000_M3 24000_28000_M3 0.018
r 24000_28000_M3 24000_32000_M3 0.018
r 24000_32000_M3 24000_36000_M3 0.018
r 24000_36000_M3 24000_40000_M3 0.018
r 24000_40000_M3 24000_44000_M3 0.018
r 24000_44000_M3 24000_48000_M3 0.018
r 24000_48000_M3 24000_52000_M3 0.018
r 24000_52000_M3 24000_56000_M3 0.018
r 24000_56000_M3 24000_60000_M3 0.018
r 24000_60000_M3 24000_64000_M3 0.018
r 24000_64000_M3 24000_68000_M3 0.018
r 24000_68000_M3 24000_72000_M3 0.018
r 24000_72000_M3 24000_76000_M3 0.018
r 24000_76000_M3 24000_80000_M3 0.018
r 24000_80000_M3 24000_84000_M3 0.018
r 24000_84000_M3 24000_88000_M3 0.018
r 24000_88000_M3 24000_92000_M3 0.018
r 24000_92000_M3 24000_96000_M3 0.018
r 24000_96000_M3 24000_100000_M3 0.018
r 28000_4000_M3 28000_8000_M3 0.018
r 28000_8000_M3 28000_12000_M3 0.018
r 28000_12000_M3 28000_16000_M3 0.018
r 28000_16000_M3 28000_20000_M3 0.018
r 28000_20000_M3 28000_24000_M3 0.018
r 28000_24000_M3 28000_28000_M3 0.018
r 28000_28000_M3 28000_32000_M3 0.018
r 28000_32000_M3 28000_36000_M3 0.018
r 28000_36000_M3 28000_40000_M3 0.018
r 28000_40000_M3 28000_44000_M3 0.018
r 28000_44000_M3 28000_48000_M3 0.018
r 28000_48000_M3 28000_52000_M3 0.018
r 28000_52000_M3 28000_56000_M3 0.018
r 28000_56000_M3 28000_60000_M3 0.018
r 28000_60000_M3 28000_64000_M3 0.018
r 28000_64000_M3 28000_68000_M3 0.018
r 28000_68000_M3 28000_72000_M3 0.018
r 28000_72000_M3 28000_76000_M3 0.018
r 28000_76000_M3 28000_80000_M3 0.018
r 28000_80000_M3 28000_84000_M3 0.018
r 28000_84000_M3 28000_88000_M3 0.018
r 28000_88000_M3 28000_92000_M3 0.018
r 28000_92000_M3 28000_96000_M3 0.018
r 28000_96000_M3 28000_100000_M3 0.018
r 32000_4000_M3 32000_8000_M3 0.018
r 32000_8000_M3 32000_12000_M3 0.018
r 32000_12000_M3 32000_16000_M3 0.018
r 32000_16000_M3 32000_20000_M3 0.018
r 32000_20000_M3 32000_24000_M3 0.018
r 32000_24000_M3 32000_28000_M3 0.018
r 32000_28000_M3 32000_32000_M3 0.018
r 32000_32000_M3 32000_36000_M3 0.018
r 32000_36000_M3 32000_40000_M3 0.018
r 32000_40000_M3 32000_44000_M3 0.018
r 32000_44000_M3 32000_48000_M3 0.018
r 32000_48000_M3 32000_52000_M3 0.018
r 32000_52000_M3 32000_56000_M3 0.018
r 32000_56000_M3 32000_60000_M3 0.018
r 32000_60000_M3 32000_64000_M3 0.018
r 32000_64000_M3 32000_68000_M3 0.018
r 32000_68000_M3 32000_72000_M3 0.018
r 32000_72000_M3 32000_76000_M3 0.018
r 32000_76000_M3 32000_80000_M3 0.018
r 32000_80000_M3 32000_84000_M3 0.018
r 32000_84000_M3 32000_88000_M3 0.018
r 32000_88000_M3 32000_92000_M3 0.018
r 32000_92000_M3 32000_96000_M3 0.018
r 32000_96000_M3 32000_100000_M3 0.018
r 36000_4000_M3 36000_8000_M3 0.018
r 36000_8000_M3 36000_12000_M3 0.018
r 36000_12000_M3 36000_16000_M3 0.018
r 36000_16000_M3 36000_20000_M3 0.018
r 36000_20000_M3 36000_24000_M3 0.018
r 36000_24000_M3 36000_28000_M3 0.018
r 36000_28000_M3 36000_32000_M3 0.018
r 36000_32000_M3 36000_36000_M3 0.018
r 36000_36000_M3 36000_40000_M3 0.018
r 36000_40000_M3 36000_44000_M3 0.018
r 36000_44000_M3 36000_48000_M3 0.018
r 36000_48000_M3 36000_52000_M3 0.018
r 36000_52000_M3 36000_56000_M3 0.018
r 36000_56000_M3 36000_60000_M3 0.018
r 36000_60000_M3 36000_64000_M3 0.018
r 36000_64000_M3 36000_68000_M3 0.018
r 36000_68000_M3 36000_72000_M3 0.018
r 36000_72000_M3 36000_76000_M3 0.018
r 36000_76000_M3 36000_80000_M3 0.018
r 36000_80000_M3 36000_84000_M3 0.018
r 36000_84000_M3 36000_88000_M3 0.018
r 36000_88000_M3 36000_92000_M3 0.018
r 36000_92000_M3 36000_96000_M3 0.018
r 36000_96000_M3 36000_100000_M3 0.018
r 40000_4000_M3 40000_8000_M3 0.018
r 40000_8000_M3 40000_12000_M3 0.018
r 40000_12000_M3 40000_16000_M3 0.018
r 40000_16000_M3 40000_20000_M3 0.018
r 40000_20000_M3 40000_24000_M3 0.018
r 40000_24000_M3 40000_28000_M3 0.018
r 40000_28000_M3 40000_32000_M3 0.018
r 40000_32000_M3 40000_36000_M3 0.018
r 40000_36000_M3 40000_40000_M3 0.018
r 40000_40000_M3 40000_44000_M3 0.018
r 40000_44000_M3 40000_48000_M3 0.018
r 40000_48000_M3 40000_52000_M3 0.018
r 40000_52000_M3 40000_56000_M3 0.018
r 40000_56000_M3 40000_60000_M3 0.018
r 40000_60000_M3 40000_64000_M3 0.018
r 40000_64000_M3 40000_68000_M3 0.018
r 40000_68000_M3 40000_72000_M3 0.018
r 40000_72000_M3 40000_76000_M3 0.018
r 40000_76000_M3 40000_80000_M3 0.018
r 40000_80000_M3 40000_84000_M3 0.018
r 40000_84000_M3 40000_88000_M3 0.018
r 40000_88000_M3 40000_92000_M3 0.018
r 40000_92000_M3 40000_96000_M3 0.018
r 40000_96000_M3 40000_100000_M3 0.018
r 44000_4000_M3 44000_8000_M3 0.018
r 44000_8000_M3 44000_12000_M3 0.018
r 44000_12000_M3 44000_16000_M3 0.018
r 44000_16000_M3 44000_20000_M3 0.018
r 44000_20000_M3 44000_24000_M3 0.018
r 44000_24000_M3 44000_28000_M3 0.018
r 44000_28000_M3 44000_32000_M3 0.018
r 44000_32000_M3 44000_36000_M3 0.018
r 44000_36000_M3 44000_40000_M3 0.018
r 44000_40000_M3 44000_44000_M3 0.018
r 44000_44000_M3 44000_48000_M3 0.018
r 44000_48000_M3 44000_52000_M3 0.018
r 44000_52000_M3 44000_56000_M3 0.018
r 44000_56000_M3 44000_60000_M3 0.018
r 44000_60000_M3 44000_64000_M3 0.018
r 44000_64000_M3 44000_68000_M3 0.018
r 44000_68000_M3 44000_72000_M3 0.018
r 44000_72000_M3 44000_76000_M3 0.018
r 44000_76000_M3 44000_80000_M3 0.018
r 44000_80000_M3 44000_84000_M3 0.018
r 44000_84000_M3 44000_88000_M3 0.018
r 44000_88000_M3 44000_92000_M3 0.018
r 44000_92000_M3 44000_96000_M3 0.018
r 44000_96000_M3 44000_100000_M3 0.018
r 48000_4000_M3 48000_8000_M3 0.018
r 48000_8000_M3 48000_12000_M3 0.018
r 48000_12000_M3 48000_16000_M3 0.018
r 48000_16000_M3 48000_20000_M3 0.018
r 48000_20000_M3 48000_24000_M3 0.018
r 48000_24000_M3 48000_28000_M3 0.018
r 48000_28000_M3 48000_32000_M3 0.018
r 48000_32000_M3 48000_36000_M3 0.018
r 48000_36000_M3 48000_40000_M3 0.018
r 48000_40000_M3 48000_44000_M3 0.018
r 48000_44000_M3 48000_48000_M3 0.018
r 48000_48000_M3 48000_52000_M3 0.018
r 48000_52000_M3 48000_56000_M3 0.018
r 48000_56000_M3 48000_60000_M3 0.018
r 48000_60000_M3 48000_64000_M3 0.018
r 48000_64000_M3 48000_68000_M3 0.018
r 48000_68000_M3 48000_72000_M3 0.018
r 48000_72000_M3 48000_76000_M3 0.018
r 48000_76000_M3 48000_80000_M3 0.018
r 48000_80000_M3 48000_84000_M3 0.018
r 48000_84000_M3 48000_88000_M3 0.018
r 48000_88000_M3 48000_92000_M3 0.018
r 48000_92000_M3 48000_96000_M3 0.018
r 48000_96000_M3 48000_100000_M3 0.018
r 52000_4000_M3 52000_8000_M3 0.018
r 52000_8000_M3 52000_12000_M3 0.018
r 52000_12000_M3 52000_16000_M3 0.018
r 52000_16000_M3 52000_20000_M3 0.018
r 52000_20000_M3 52000_24000_M3 0.018
r 52000_24000_M3 52000_28000_M3 0.018
r 52000_28000_M3 52000_32000_M3 0.018
r 52000_32000_M3 52000_36000_M3 0.018
r 52000_36000_M3 52000_40000_M3 0.018
r 52000_40000_M3 52000_44000_M3 0.018
r 52000_44000_M3 52000_48000_M3 0.018
r 52000_48000_M3 52000_52000_M3 0.018
r 52000_52000_M3 52000_56000_M3 0.018
r 52000_56000_M3 52000_60000_M3 0.018
r 52000_60000_M3 52000_64000_M3 0.018
r 52000_64000_M3 52000_68000_M3 0.018
r 52000_68000_M3 52000_72000_M3 0.018
r 52000_72000_M3 52000_76000_M3 0.018
r 52000_76000_M3 52000_80000_M3 0.018
r 52000_80000_M3 52000_84000_M3 0.018
r 52000_84000_M3 52000_88000_M3 0.018
r 52000_88000_M3 52000_92000_M3 0.018
r 52000_92000_M3 52000_96000_M3 0.018
r 52000_96000_M3 52000_100000_M3 0.018
r 56000_4000_M3 56000_8000_M3 0.018
r 56000_8000_M3 56000_12000_M3 0.018
r 56000_12000_M3 56000_16000_M3 0.018
r 56000_16000_M3 56000_20000_M3 0.018
r 56000_20000_M3 56000_24000_M3 0.018
r 56000_24000_M3 56000_28000_M3 0.018
r 56000_28000_M3 56000_32000_M3 0.018
r 56000_32000_M3 56000_36000_M3 0.018
r 56000_36000_M3 56000_40000_M3 0.018
r 56000_40000_M3 56000_44000_M3 0.018
r 56000_44000_M3 56000_48000_M3 0.018
r 56000_48000_M3 56000_52000_M3 0.018
r 56000_52000_M3 56000_56000_M3 0.018
r 56000_56000_M3 56000_60000_M3 0.018
r 56000_60000_M3 56000_64000_M3 0.018
r 56000_64000_M3 56000_68000_M3 0.018
r 56000_68000_M3 56000_72000_M3 0.018
r 56000_72000_M3 56000_76000_M3 0.018
r 56000_76000_M3 56000_80000_M3 0.018
r 56000_80000_M3 56000_84000_M3 0.018
r 56000_84000_M3 56000_88000_M3 0.018
r 56000_88000_M3 56000_92000_M3 0.018
r 56000_92000_M3 56000_96000_M3 0.018
r 56000_96000_M3 56000_100000_M3 0.018
r 60000_4000_M3 60000_8000_M3 0.018
r 60000_8000_M3 60000_12000_M3 0.018
r 60000_12000_M3 60000_16000_M3 0.018
r 60000_16000_M3 60000_20000_M3 0.018
r 60000_20000_M3 60000_24000_M3 0.018
r 60000_24000_M3 60000_28000_M3 0.018
r 60000_28000_M3 60000_32000_M3 0.018
r 60000_32000_M3 60000_36000_M3 0.018
r 60000_36000_M3 60000_40000_M3 0.018
r 60000_40000_M3 60000_44000_M3 0.018
r 60000_44000_M3 60000_48000_M3 0.018
r 60000_48000_M3 60000_52000_M3 0.018
r 60000_52000_M3 60000_56000_M3 0.018
r 60000_56000_M3 60000_60000_M3 0.018
r 60000_60000_M3 60000_64000_M3 0.018
r 60000_64000_M3 60000_68000_M3 0.018
r 60000_68000_M3 60000_72000_M3 0.018
r 60000_72000_M3 60000_76000_M3 0.018
r 60000_76000_M3 60000_80000_M3 0.018
r 60000_80000_M3 60000_84000_M3 0.018
r 60000_84000_M3 60000_88000_M3 0.018
r 60000_88000_M3 60000_92000_M3 0.018
r 60000_92000_M3 60000_96000_M3 0.018
r 60000_96000_M3 60000_100000_M3 0.018
r 64000_4000_M3 64000_8000_M3 0.018
r 64000_8000_M3 64000_12000_M3 0.018
r 64000_12000_M3 64000_16000_M3 0.018
r 64000_16000_M3 64000_20000_M3 0.018
r 64000_20000_M3 64000_24000_M3 0.018
r 64000_24000_M3 64000_28000_M3 0.018
r 64000_28000_M3 64000_32000_M3 0.018
r 64000_32000_M3 64000_36000_M3 0.018
r 64000_36000_M3 64000_40000_M3 0.018
r 64000_40000_M3 64000_44000_M3 0.018
r 64000_44000_M3 64000_48000_M3 0.018
r 64000_48000_M3 64000_52000_M3 0.018
r 64000_52000_M3 64000_56000_M3 0.018
r 64000_56000_M3 64000_60000_M3 0.018
r 64000_60000_M3 64000_64000_M3 0.018
r 64000_64000_M3 64000_68000_M3 0.018
r 64000_68000_M3 64000_72000_M3 0.018
r 64000_72000_M3 64000_76000_M3 0.018
r 64000_76000_M3 64000_80000_M3 0.018
r 64000_80000_M3 64000_84000_M3 0.018
r 64000_84000_M3 64000_88000_M3 0.018
r 64000_88000_M3 64000_92000_M3 0.018
r 64000_92000_M3 64000_96000_M3 0.018
r 64000_96000_M3 64000_100000_M3 0.018
r 68000_4000_M3 68000_8000_M3 0.018
r 68000_8000_M3 68000_12000_M3 0.018
r 68000_12000_M3 68000_16000_M3 0.018
r 68000_16000_M3 68000_20000_M3 0.018
r 68000_20000_M3 68000_24000_M3 0.018
r 68000_24000_M3 68000_28000_M3 0.018
r 68000_28000_M3 68000_32000_M3 0.018
r 68000_32000_M3 68000_36000_M3 0.018
r 68000_36000_M3 68000_40000_M3 0.018
r 68000_40000_M3 68000_44000_M3 0.018
r 68000_44000_M3 68000_48000_M3 0.018
r 68000_48000_M3 68000_52000_M3 0.018
r 68000_52000_M3 68000_56000_M3 0.018
r 68000_56000_M3 68000_60000_M3 0.018
r 68000_60000_M3 68000_64000_M3 0.018
r 68000_64000_M3 68000_68000_M3 0.018
r 68000_68000_M3 68000_72000_M3 0.018
r 68000_72000_M3 68000_76000_M3 0.018
r 68000_76000_M3 68000_80000_M3 0.018
r 68000_80000_M3 68000_84000_M3 0.018
r 68000_84000_M3 68000_88000_M3 0.018
r 68000_88000_M3 68000_92000_M3 0.018
r 68000_92000_M3 68000_96000_M3 0.018
r 68000_96000_M3 68000_100000_M3 0.018
r 72000_4000_M3 72000_8000_M3 0.018
r 72000_8000_M3 72000_12000_M3 0.018
r 72000_12000_M3 72000_16000_M3 0.018
r 72000_16000_M3 72000_20000_M3 0.018
r 72000_20000_M3 72000_24000_M3 0.018
r 72000_24000_M3 72000_28000_M3 0.018
r 72000_28000_M3 72000_32000_M3 0.018
r 72000_32000_M3 72000_36000_M3 0.018
r 72000_36000_M3 72000_40000_M3 0.018
r 72000_40000_M3 72000_44000_M3 0.018
r 72000_44000_M3 72000_48000_M3 0.018
r 72000_48000_M3 72000_52000_M3 0.018
r 72000_52000_M3 72000_56000_M3 0.018
r 72000_56000_M3 72000_60000_M3 0.018
r 72000_60000_M3 72000_64000_M3 0.018
r 72000_64000_M3 72000_68000_M3 0.018
r 72000_68000_M3 72000_72000_M3 0.018
r 72000_72000_M3 72000_76000_M3 0.018
r 72000_76000_M3 72000_80000_M3 0.018
r 72000_80000_M3 72000_84000_M3 0.018
r 72000_84000_M3 72000_88000_M3 0.018
r 72000_88000_M3 72000_92000_M3 0.018
r 72000_92000_M3 72000_96000_M3 0.018
r 72000_96000_M3 72000_100000_M3 0.018
r 76000_4000_M3 76000_8000_M3 0.018
r 76000_8000_M3 76000_12000_M3 0.018
r 76000_12000_M3 76000_16000_M3 0.018
r 76000_16000_M3 76000_20000_M3 0.018
r 76000_20000_M3 76000_24000_M3 0.018
r 76000_24000_M3 76000_28000_M3 0.018
r 76000_28000_M3 76000_32000_M3 0.018
r 76000_32000_M3 76000_36000_M3 0.018
r 76000_36000_M3 76000_40000_M3 0.018
r 76000_40000_M3 76000_44000_M3 0.018
r 76000_44000_M3 76000_48000_M3 0.018
r 76000_48000_M3 76000_52000_M3 0.018
r 76000_52000_M3 76000_56000_M3 0.018
r 76000_56000_M3 76000_60000_M3 0.018
r 76000_60000_M3 76000_64000_M3 0.018
r 76000_64000_M3 76000_68000_M3 0.018
r 76000_68000_M3 76000_72000_M3 0.018
r 76000_72000_M3 76000_76000_M3 0.018
r 76000_76000_M3 76000_80000_M3 0.018
r 76000_80000_M3 76000_84000_M3 0.018
r 76000_84000_M3 76000_88000_M3 0.018
r 76000_88000_M3 76000_92000_M3 0.018
r 76000_92000_M3 76000_96000_M3 0.018
r 76000_96000_M3 76000_100000_M3 0.018
r 80000_4000_M3 80000_8000_M3 0.018
r 80000_8000_M3 80000_12000_M3 0.018
r 80000_12000_M3 80000_16000_M3 0.018
r 80000_16000_M3 80000_20000_M3 0.018
r 80000_20000_M3 80000_24000_M3 0.018
r 80000_24000_M3 80000_28000_M3 0.018
r 80000_28000_M3 80000_32000_M3 0.018
r 80000_32000_M3 80000_36000_M3 0.018
r 80000_36000_M3 80000_40000_M3 0.018
r 80000_40000_M3 80000_44000_M3 0.018
r 80000_44000_M3 80000_48000_M3 0.018
r 80000_48000_M3 80000_52000_M3 0.018
r 80000_52000_M3 80000_56000_M3 0.018
r 80000_56000_M3 80000_60000_M3 0.018
r 80000_60000_M3 80000_64000_M3 0.018
r 80000_64000_M3 80000_68000_M3 0.018
r 80000_68000_M3 80000_72000_M3 0.018
r 80000_72000_M3 80000_76000_M3 0.018
r 80000_76000_M3 80000_80000_M3 0.018
r 80000_80000_M3 80000_84000_M3 0.018
r 80000_84000_M3 80000_88000_M3 0.018
r 80000_88000_M3 80000_92000_M3 0.018
r 80000_92000_M3 80000_96000_M3 0.018
r 80000_96000_M3 80000_100000_M3 0.018
r 84000_4000_M3 84000_8000_M3 0.018
r 84000_8000_M3 84000_12000_M3 0.018
r 84000_12000_M3 84000_16000_M3 0.018
r 84000_16000_M3 84000_20000_M3 0.018
r 84000_20000_M3 84000_24000_M3 0.018
r 84000_24000_M3 84000_28000_M3 0.018
r 84000_28000_M3 84000_32000_M3 0.018
r 84000_32000_M3 84000_36000_M3 0.018
r 84000_36000_M3 84000_40000_M3 0.018
r 84000_40000_M3 84000_44000_M3 0.018
r 84000_44000_M3 84000_48000_M3 0.018
r 84000_48000_M3 84000_52000_M3 0.018
r 84000_52000_M3 84000_56000_M3 0.018
r 84000_56000_M3 84000_60000_M3 0.018
r 84000_60000_M3 84000_64000_M3 0.018
r 84000_64000_M3 84000_68000_M3 0.018
r 84000_68000_M3 84000_72000_M3 0.018
r 84000_72000_M3 84000_76000_M3 0.018
r 84000_76000_M3 84000_80000_M3 0.018
r 84000_80000_M3 84000_84000_M3 0.018
r 84000_84000_M3 84000_88000_M3 0.018
r 84000_88000_M3 84000_92000_M3 0.018
r 84000_92000_M3 84000_96000_M3 0.018
r 84000_96000_M3 84000_100000_M3 0.018
r 88000_4000_M3 88000_8000_M3 0.018
r 88000_8000_M3 88000_12000_M3 0.018
r 88000_12000_M3 88000_16000_M3 0.018
r 88000_16000_M3 88000_20000_M3 0.018
r 88000_20000_M3 88000_24000_M3 0.018
r 88000_24000_M3 88000_28000_M3 0.018
r 88000_28000_M3 88000_32000_M3 0.018
r 88000_32000_M3 88000_36000_M3 0.018
r 88000_36000_M3 88000_40000_M3 0.018
r 88000_40000_M3 88000_44000_M3 0.018
r 88000_44000_M3 88000_48000_M3 0.018
r 88000_48000_M3 88000_52000_M3 0.018
r 88000_52000_M3 88000_56000_M3 0.018
r 88000_56000_M3 88000_60000_M3 0.018
r 88000_60000_M3 88000_64000_M3 0.018
r 88000_64000_M3 88000_68000_M3 0.018
r 88000_68000_M3 88000_72000_M3 0.018
r 88000_72000_M3 88000_76000_M3 0.018
r 88000_76000_M3 88000_80000_M3 0.018
r 88000_80000_M3 88000_84000_M3 0.018
r 88000_84000_M3 88000_88000_M3 0.018
r 88000_88000_M3 88000_92000_M3 0.018
r 88000_92000_M3 88000_96000_M3 0.018
r 88000_96000_M3 88000_100000_M3 0.018
r 92000_4000_M3 92000_8000_M3 0.018
r 92000_8000_M3 92000_12000_M3 0.018
r 92000_12000_M3 92000_16000_M3 0.018
r 92000_16000_M3 92000_20000_M3 0.018
r 92000_20000_M3 92000_24000_M3 0.018
r 92000_24000_M3 92000_28000_M3 0.018
r 92000_28000_M3 92000_32000_M3 0.018
r 92000_32000_M3 92000_36000_M3 0.018
r 92000_36000_M3 92000_40000_M3 0.018
r 92000_40000_M3 92000_44000_M3 0.018
r 92000_44000_M3 92000_48000_M3 0.018
r 92000_48000_M3 92000_52000_M3 0.018
r 92000_52000_M3 92000_56000_M3 0.018
r 92000_56000_M3 92000_60000_M3 0.018
r 92000_60000_M3 92000_64000_M3 0.018
r 92000_64000_M3 92000_68000_M3 0.018
r 92000_68000_M3 92000_72000_M3 0.018
r 92000_72000_M3 92000_76000_M3 0.018
r 92000_76000_M3 92000_80000_M3 0.018
r 92000_80000_M3 92000_84000_M3 0.018
r 92000_84000_M3 92000_88000_M3 0.018
r 92000_88000_M3 92000_92000_M3 0.018
r 92000_92000_M3 92000_96000_M3 0.018
r 92000_96000_M3 92000_100000_M3 0.018
r 96000_4000_M3 96000_8000_M3 0.018
r 96000_8000_M3 96000_12000_M3 0.018
r 96000_12000_M3 96000_16000_M3 0.018
r 96000_16000_M3 96000_20000_M3 0.018
r 96000_20000_M3 96000_24000_M3 0.018
r 96000_24000_M3 96000_28000_M3 0.018
r 96000_28000_M3 96000_32000_M3 0.018
r 96000_32000_M3 96000_36000_M3 0.018
r 96000_36000_M3 96000_40000_M3 0.018
r 96000_40000_M3 96000_44000_M3 0.018
r 96000_44000_M3 96000_48000_M3 0.018
r 96000_48000_M3 96000_52000_M3 0.018
r 96000_52000_M3 96000_56000_M3 0.018
r 96000_56000_M3 96000_60000_M3 0.018
r 96000_60000_M3 96000_64000_M3 0.018
r 96000_64000_M3 96000_68000_M3 0.018
r 96000_68000_M3 96000_72000_M3 0.018
r 96000_72000_M3 96000_76000_M3 0.018
r 96000_76000_M3 96000_80000_M3 0.018
r 96000_80000_M3 96000_84000_M3 0.018
r 96000_84000_M3 96000_88000_M3 0.018
r 96000_88000_M3 96000_92000_M3 0.018
r 96000_92000_M3 96000_96000_M3 0.018
r 96000_96000_M3 96000_100000_M3 0.018
r 100000_4000_M3 100000_8000_M3 0.018
r 100000_8000_M3 100000_12000_M3 0.018
r 100000_12000_M3 100000_16000_M3 0.018
r 100000_16000_M3 100000_20000_M3 0.018
r 100000_20000_M3 100000_24000_M3 0.018
r 100000_24000_M3 100000_28000_M3 0.018
r 100000_28000_M3 100000_32000_M3 0.018
r 100000_32000_M3 100000_36000_M3 0.018
r 100000_36000_M3 100000_40000_M3 0.018
r 100000_40000_M3 100000_44000_M3 0.018
r 100000_44000_M3 100000_48000_M3 0.018
r 100000_48000_M3 100000_52000_M3 0.018
r 100000_52000_M3 100000_56000_M3 0.018
r 100000_56000_M3 100000_60000_M3 0.018
r 100000_60000_M3 100000_64000_M3 0.018
r 100000_64000_M3 100000_68000_M3 0.018
r 100000_68000_M3 100000_72000_M3 0.018
r 100000_72000_M3 100000_76000_M3 0.018
r 100000_76000_M3 100000_80000_M3 0.018
r 100000_80000_M3 100000_84000_M3 0.018
r 100000_84000_M3 100000_88000_M3 0.018
r 100000_88000_M3 100000_92000_M3 0.018
r 100000_92000_M3 100000_96000_M3 0.018
r 100000_96000_M3 100000_100000_M3 0.018

* ============================================================================
* Layer M4 - 25x25 grid
* ============================================================================

* M4 Horizontal resistors
r 4000_4000_M4 8000_4000_M4 0.012
r 8000_4000_M4 12000_4000_M4 0.012
r 12000_4000_M4 16000_4000_M4 0.012
r 16000_4000_M4 20000_4000_M4 0.012
r 20000_4000_M4 24000_4000_M4 0.012
r 24000_4000_M4 28000_4000_M4 0.012
r 28000_4000_M4 32000_4000_M4 0.012
r 32000_4000_M4 36000_4000_M4 0.012
r 36000_4000_M4 40000_4000_M4 0.012
r 40000_4000_M4 44000_4000_M4 0.012
r 44000_4000_M4 48000_4000_M4 0.012
r 48000_4000_M4 52000_4000_M4 0.012
r 52000_4000_M4 56000_4000_M4 0.012
r 56000_4000_M4 60000_4000_M4 0.012
r 60000_4000_M4 64000_4000_M4 0.012
r 64000_4000_M4 68000_4000_M4 0.012
r 68000_4000_M4 72000_4000_M4 0.012
r 72000_4000_M4 76000_4000_M4 0.012
r 76000_4000_M4 80000_4000_M4 0.012
r 80000_4000_M4 84000_4000_M4 0.012
r 84000_4000_M4 88000_4000_M4 0.012
r 88000_4000_M4 92000_4000_M4 0.012
r 92000_4000_M4 96000_4000_M4 0.012
r 96000_4000_M4 100000_4000_M4 0.012
r 4000_8000_M4 8000_8000_M4 0.012
r 8000_8000_M4 12000_8000_M4 0.012
r 12000_8000_M4 16000_8000_M4 0.012
r 16000_8000_M4 20000_8000_M4 0.012
r 20000_8000_M4 24000_8000_M4 0.012
r 24000_8000_M4 28000_8000_M4 0.012
r 28000_8000_M4 32000_8000_M4 0.012
r 32000_8000_M4 36000_8000_M4 0.012
r 36000_8000_M4 40000_8000_M4 0.012
r 40000_8000_M4 44000_8000_M4 0.012
r 44000_8000_M4 48000_8000_M4 0.012
r 48000_8000_M4 52000_8000_M4 0.012
r 52000_8000_M4 56000_8000_M4 0.012
r 56000_8000_M4 60000_8000_M4 0.012
r 60000_8000_M4 64000_8000_M4 0.012
r 64000_8000_M4 68000_8000_M4 0.012
r 68000_8000_M4 72000_8000_M4 0.012
r 72000_8000_M4 76000_8000_M4 0.012
r 76000_8000_M4 80000_8000_M4 0.012
r 80000_8000_M4 84000_8000_M4 0.012
r 84000_8000_M4 88000_8000_M4 0.012
r 88000_8000_M4 92000_8000_M4 0.012
r 92000_8000_M4 96000_8000_M4 0.012
r 96000_8000_M4 100000_8000_M4 0.012
r 4000_12000_M4 8000_12000_M4 0.012
r 8000_12000_M4 12000_12000_M4 0.012
r 12000_12000_M4 16000_12000_M4 0.012
r 16000_12000_M4 20000_12000_M4 0.012
r 20000_12000_M4 24000_12000_M4 0.012
r 24000_12000_M4 28000_12000_M4 0.012
r 28000_12000_M4 32000_12000_M4 0.012
r 32000_12000_M4 36000_12000_M4 0.012
r 36000_12000_M4 40000_12000_M4 0.012
r 40000_12000_M4 44000_12000_M4 0.012
r 44000_12000_M4 48000_12000_M4 0.012
r 48000_12000_M4 52000_12000_M4 0.012
r 52000_12000_M4 56000_12000_M4 0.012
r 56000_12000_M4 60000_12000_M4 0.012
r 60000_12000_M4 64000_12000_M4 0.012
r 64000_12000_M4 68000_12000_M4 0.012
r 68000_12000_M4 72000_12000_M4 0.012
r 72000_12000_M4 76000_12000_M4 0.012
r 76000_12000_M4 80000_12000_M4 0.012
r 80000_12000_M4 84000_12000_M4 0.012
r 84000_12000_M4 88000_12000_M4 0.012
r 88000_12000_M4 92000_12000_M4 0.012
r 92000_12000_M4 96000_12000_M4 0.012
r 96000_12000_M4 100000_12000_M4 0.012
r 4000_16000_M4 8000_16000_M4 0.012
r 8000_16000_M4 12000_16000_M4 0.012
r 12000_16000_M4 16000_16000_M4 0.012
r 16000_16000_M4 20000_16000_M4 0.012
r 20000_16000_M4 24000_16000_M4 0.012
r 24000_16000_M4 28000_16000_M4 0.012
r 28000_16000_M4 32000_16000_M4 0.012
r 32000_16000_M4 36000_16000_M4 0.012
r 36000_16000_M4 40000_16000_M4 0.012
r 40000_16000_M4 44000_16000_M4 0.012
r 44000_16000_M4 48000_16000_M4 0.012
r 48000_16000_M4 52000_16000_M4 0.012
r 52000_16000_M4 56000_16000_M4 0.012
r 56000_16000_M4 60000_16000_M4 0.012
r 60000_16000_M4 64000_16000_M4 0.012
r 64000_16000_M4 68000_16000_M4 0.012
r 68000_16000_M4 72000_16000_M4 0.012
r 72000_16000_M4 76000_16000_M4 0.012
r 76000_16000_M4 80000_16000_M4 0.012
r 80000_16000_M4 84000_16000_M4 0.012
r 84000_16000_M4 88000_16000_M4 0.012
r 88000_16000_M4 92000_16000_M4 0.012
r 92000_16000_M4 96000_16000_M4 0.012
r 96000_16000_M4 100000_16000_M4 0.012
r 4000_20000_M4 8000_20000_M4 0.012
r 8000_20000_M4 12000_20000_M4 0.012
r 12000_20000_M4 16000_20000_M4 0.012
r 16000_20000_M4 20000_20000_M4 0.012
r 20000_20000_M4 24000_20000_M4 0.012
r 24000_20000_M4 28000_20000_M4 0.012
r 28000_20000_M4 32000_20000_M4 0.012
r 32000_20000_M4 36000_20000_M4 0.012
r 36000_20000_M4 40000_20000_M4 0.012
r 40000_20000_M4 44000_20000_M4 0.012
r 44000_20000_M4 48000_20000_M4 0.012
r 48000_20000_M4 52000_20000_M4 0.012
r 52000_20000_M4 56000_20000_M4 0.012
r 56000_20000_M4 60000_20000_M4 0.012
r 60000_20000_M4 64000_20000_M4 0.012
r 64000_20000_M4 68000_20000_M4 0.012
r 68000_20000_M4 72000_20000_M4 0.012
r 72000_20000_M4 76000_20000_M4 0.012
r 76000_20000_M4 80000_20000_M4 0.012
r 80000_20000_M4 84000_20000_M4 0.012
r 84000_20000_M4 88000_20000_M4 0.012
r 88000_20000_M4 92000_20000_M4 0.012
r 92000_20000_M4 96000_20000_M4 0.012
r 96000_20000_M4 100000_20000_M4 0.012
r 4000_24000_M4 8000_24000_M4 0.012
r 8000_24000_M4 12000_24000_M4 0.012
r 12000_24000_M4 16000_24000_M4 0.012
r 16000_24000_M4 20000_24000_M4 0.012
r 20000_24000_M4 24000_24000_M4 0.012
r 24000_24000_M4 28000_24000_M4 0.012
r 28000_24000_M4 32000_24000_M4 0.012
r 32000_24000_M4 36000_24000_M4 0.012
r 36000_24000_M4 40000_24000_M4 0.012
r 40000_24000_M4 44000_24000_M4 0.012
r 44000_24000_M4 48000_24000_M4 0.012
r 48000_24000_M4 52000_24000_M4 0.012
r 52000_24000_M4 56000_24000_M4 0.012
r 56000_24000_M4 60000_24000_M4 0.012
r 60000_24000_M4 64000_24000_M4 0.012
r 64000_24000_M4 68000_24000_M4 0.012
r 68000_24000_M4 72000_24000_M4 0.012
r 72000_24000_M4 76000_24000_M4 0.012
r 76000_24000_M4 80000_24000_M4 0.012
r 80000_24000_M4 84000_24000_M4 0.012
r 84000_24000_M4 88000_24000_M4 0.012
r 88000_24000_M4 92000_24000_M4 0.012
r 92000_24000_M4 96000_24000_M4 0.012
r 96000_24000_M4 100000_24000_M4 0.012
r 4000_28000_M4 8000_28000_M4 0.012
r 8000_28000_M4 12000_28000_M4 0.012
r 12000_28000_M4 16000_28000_M4 0.012
r 16000_28000_M4 20000_28000_M4 0.012
r 20000_28000_M4 24000_28000_M4 0.012
r 24000_28000_M4 28000_28000_M4 0.012
r 28000_28000_M4 32000_28000_M4 0.012
r 32000_28000_M4 36000_28000_M4 0.012
r 36000_28000_M4 40000_28000_M4 0.012
r 40000_28000_M4 44000_28000_M4 0.012
r 44000_28000_M4 48000_28000_M4 0.012
r 48000_28000_M4 52000_28000_M4 0.012
r 52000_28000_M4 56000_28000_M4 0.012
r 56000_28000_M4 60000_28000_M4 0.012
r 60000_28000_M4 64000_28000_M4 0.012
r 64000_28000_M4 68000_28000_M4 0.012
r 68000_28000_M4 72000_28000_M4 0.012
r 72000_28000_M4 76000_28000_M4 0.012
r 76000_28000_M4 80000_28000_M4 0.012
r 80000_28000_M4 84000_28000_M4 0.012
r 84000_28000_M4 88000_28000_M4 0.012
r 88000_28000_M4 92000_28000_M4 0.012
r 92000_28000_M4 96000_28000_M4 0.012
r 96000_28000_M4 100000_28000_M4 0.012
r 4000_32000_M4 8000_32000_M4 0.012
r 8000_32000_M4 12000_32000_M4 0.012
r 12000_32000_M4 16000_32000_M4 0.012
r 16000_32000_M4 20000_32000_M4 0.012
r 20000_32000_M4 24000_32000_M4 0.012
r 24000_32000_M4 28000_32000_M4 0.012
r 28000_32000_M4 32000_32000_M4 0.012
r 32000_32000_M4 36000_32000_M4 0.012
r 36000_32000_M4 40000_32000_M4 0.012
r 40000_32000_M4 44000_32000_M4 0.012
r 44000_32000_M4 48000_32000_M4 0.012
r 48000_32000_M4 52000_32000_M4 0.012
r 52000_32000_M4 56000_32000_M4 0.012
r 56000_32000_M4 60000_32000_M4 0.012
r 60000_32000_M4 64000_32000_M4 0.012
r 64000_32000_M4 68000_32000_M4 0.012
r 68000_32000_M4 72000_32000_M4 0.012
r 72000_32000_M4 76000_32000_M4 0.012
r 76000_32000_M4 80000_32000_M4 0.012
r 80000_32000_M4 84000_32000_M4 0.012
r 84000_32000_M4 88000_32000_M4 0.012
r 88000_32000_M4 92000_32000_M4 0.012
r 92000_32000_M4 96000_32000_M4 0.012
r 96000_32000_M4 100000_32000_M4 0.012
r 4000_36000_M4 8000_36000_M4 0.012
r 8000_36000_M4 12000_36000_M4 0.012
r 12000_36000_M4 16000_36000_M4 0.012
r 16000_36000_M4 20000_36000_M4 0.012
r 20000_36000_M4 24000_36000_M4 0.012
r 24000_36000_M4 28000_36000_M4 0.012
r 28000_36000_M4 32000_36000_M4 0.012
r 32000_36000_M4 36000_36000_M4 0.012
r 36000_36000_M4 40000_36000_M4 0.012
r 40000_36000_M4 44000_36000_M4 0.012
r 44000_36000_M4 48000_36000_M4 0.012
r 48000_36000_M4 52000_36000_M4 0.012
r 52000_36000_M4 56000_36000_M4 0.012
r 56000_36000_M4 60000_36000_M4 0.012
r 60000_36000_M4 64000_36000_M4 0.012
r 64000_36000_M4 68000_36000_M4 0.012
r 68000_36000_M4 72000_36000_M4 0.012
r 72000_36000_M4 76000_36000_M4 0.012
r 76000_36000_M4 80000_36000_M4 0.012
r 80000_36000_M4 84000_36000_M4 0.012
r 84000_36000_M4 88000_36000_M4 0.012
r 88000_36000_M4 92000_36000_M4 0.012
r 92000_36000_M4 96000_36000_M4 0.012
r 96000_36000_M4 100000_36000_M4 0.012
r 4000_40000_M4 8000_40000_M4 0.012
r 8000_40000_M4 12000_40000_M4 0.012
r 12000_40000_M4 16000_40000_M4 0.012
r 16000_40000_M4 20000_40000_M4 0.012
r 20000_40000_M4 24000_40000_M4 0.012
r 24000_40000_M4 28000_40000_M4 0.012
r 28000_40000_M4 32000_40000_M4 0.012
r 32000_40000_M4 36000_40000_M4 0.012
r 36000_40000_M4 40000_40000_M4 0.012
r 40000_40000_M4 44000_40000_M4 0.012
r 44000_40000_M4 48000_40000_M4 0.012
r 48000_40000_M4 52000_40000_M4 0.012
r 52000_40000_M4 56000_40000_M4 0.012
r 56000_40000_M4 60000_40000_M4 0.012
r 60000_40000_M4 64000_40000_M4 0.012
r 64000_40000_M4 68000_40000_M4 0.012
r 68000_40000_M4 72000_40000_M4 0.012
r 72000_40000_M4 76000_40000_M4 0.012
r 76000_40000_M4 80000_40000_M4 0.012
r 80000_40000_M4 84000_40000_M4 0.012
r 84000_40000_M4 88000_40000_M4 0.012
r 88000_40000_M4 92000_40000_M4 0.012
r 92000_40000_M4 96000_40000_M4 0.012
r 96000_40000_M4 100000_40000_M4 0.012
r 4000_44000_M4 8000_44000_M4 0.012
r 8000_44000_M4 12000_44000_M4 0.012
r 12000_44000_M4 16000_44000_M4 0.012
r 16000_44000_M4 20000_44000_M4 0.012
r 20000_44000_M4 24000_44000_M4 0.012
r 24000_44000_M4 28000_44000_M4 0.012
r 28000_44000_M4 32000_44000_M4 0.012
r 32000_44000_M4 36000_44000_M4 0.012
r 36000_44000_M4 40000_44000_M4 0.012
r 40000_44000_M4 44000_44000_M4 0.012
r 44000_44000_M4 48000_44000_M4 0.012
r 48000_44000_M4 52000_44000_M4 0.012
r 52000_44000_M4 56000_44000_M4 0.012
r 56000_44000_M4 60000_44000_M4 0.012
r 60000_44000_M4 64000_44000_M4 0.012
r 64000_44000_M4 68000_44000_M4 0.012
r 68000_44000_M4 72000_44000_M4 0.012
r 72000_44000_M4 76000_44000_M4 0.012
r 76000_44000_M4 80000_44000_M4 0.012
r 80000_44000_M4 84000_44000_M4 0.012
r 84000_44000_M4 88000_44000_M4 0.012
r 88000_44000_M4 92000_44000_M4 0.012
r 92000_44000_M4 96000_44000_M4 0.012
r 96000_44000_M4 100000_44000_M4 0.012
r 4000_48000_M4 8000_48000_M4 0.012
r 8000_48000_M4 12000_48000_M4 0.012
r 12000_48000_M4 16000_48000_M4 0.012
r 16000_48000_M4 20000_48000_M4 0.012
r 20000_48000_M4 24000_48000_M4 0.012
r 24000_48000_M4 28000_48000_M4 0.012
r 28000_48000_M4 32000_48000_M4 0.012
r 32000_48000_M4 36000_48000_M4 0.012
r 36000_48000_M4 40000_48000_M4 0.012
r 40000_48000_M4 44000_48000_M4 0.012
r 44000_48000_M4 48000_48000_M4 0.012
r 48000_48000_M4 52000_48000_M4 0.012
r 52000_48000_M4 56000_48000_M4 0.012
r 56000_48000_M4 60000_48000_M4 0.012
r 60000_48000_M4 64000_48000_M4 0.012
r 64000_48000_M4 68000_48000_M4 0.012
r 68000_48000_M4 72000_48000_M4 0.012
r 72000_48000_M4 76000_48000_M4 0.012
r 76000_48000_M4 80000_48000_M4 0.012
r 80000_48000_M4 84000_48000_M4 0.012
r 84000_48000_M4 88000_48000_M4 0.012
r 88000_48000_M4 92000_48000_M4 0.012
r 92000_48000_M4 96000_48000_M4 0.012
r 96000_48000_M4 100000_48000_M4 0.012
r 4000_52000_M4 8000_52000_M4 0.012
r 8000_52000_M4 12000_52000_M4 0.012
r 12000_52000_M4 16000_52000_M4 0.012
r 16000_52000_M4 20000_52000_M4 0.012
r 20000_52000_M4 24000_52000_M4 0.012
r 24000_52000_M4 28000_52000_M4 0.012
r 28000_52000_M4 32000_52000_M4 0.012
r 32000_52000_M4 36000_52000_M4 0.012
r 36000_52000_M4 40000_52000_M4 0.012
r 40000_52000_M4 44000_52000_M4 0.012
r 44000_52000_M4 48000_52000_M4 0.012
r 48000_52000_M4 52000_52000_M4 0.012
r 52000_52000_M4 56000_52000_M4 0.012
r 56000_52000_M4 60000_52000_M4 0.012
r 60000_52000_M4 64000_52000_M4 0.012
r 64000_52000_M4 68000_52000_M4 0.012
r 68000_52000_M4 72000_52000_M4 0.012
r 72000_52000_M4 76000_52000_M4 0.012
r 76000_52000_M4 80000_52000_M4 0.012
r 80000_52000_M4 84000_52000_M4 0.012
r 84000_52000_M4 88000_52000_M4 0.012
r 88000_52000_M4 92000_52000_M4 0.012
r 92000_52000_M4 96000_52000_M4 0.012
r 96000_52000_M4 100000_52000_M4 0.012
r 4000_56000_M4 8000_56000_M4 0.012
r 8000_56000_M4 12000_56000_M4 0.012
r 12000_56000_M4 16000_56000_M4 0.012
r 16000_56000_M4 20000_56000_M4 0.012
r 20000_56000_M4 24000_56000_M4 0.012
r 24000_56000_M4 28000_56000_M4 0.012
r 28000_56000_M4 32000_56000_M4 0.012
r 32000_56000_M4 36000_56000_M4 0.012
r 36000_56000_M4 40000_56000_M4 0.012
r 40000_56000_M4 44000_56000_M4 0.012
r 44000_56000_M4 48000_56000_M4 0.012
r 48000_56000_M4 52000_56000_M4 0.012
r 52000_56000_M4 56000_56000_M4 0.012
r 56000_56000_M4 60000_56000_M4 0.012
r 60000_56000_M4 64000_56000_M4 0.012
r 64000_56000_M4 68000_56000_M4 0.012
r 68000_56000_M4 72000_56000_M4 0.012
r 72000_56000_M4 76000_56000_M4 0.012
r 76000_56000_M4 80000_56000_M4 0.012
r 80000_56000_M4 84000_56000_M4 0.012
r 84000_56000_M4 88000_56000_M4 0.012
r 88000_56000_M4 92000_56000_M4 0.012
r 92000_56000_M4 96000_56000_M4 0.012
r 96000_56000_M4 100000_56000_M4 0.012
r 4000_60000_M4 8000_60000_M4 0.012
r 8000_60000_M4 12000_60000_M4 0.012
r 12000_60000_M4 16000_60000_M4 0.012
r 16000_60000_M4 20000_60000_M4 0.012
r 20000_60000_M4 24000_60000_M4 0.012
r 24000_60000_M4 28000_60000_M4 0.012
r 28000_60000_M4 32000_60000_M4 0.012
r 32000_60000_M4 36000_60000_M4 0.012
r 36000_60000_M4 40000_60000_M4 0.012
r 40000_60000_M4 44000_60000_M4 0.012
r 44000_60000_M4 48000_60000_M4 0.012
r 48000_60000_M4 52000_60000_M4 0.012
r 52000_60000_M4 56000_60000_M4 0.012
r 56000_60000_M4 60000_60000_M4 0.012
r 60000_60000_M4 64000_60000_M4 0.012
r 64000_60000_M4 68000_60000_M4 0.012
r 68000_60000_M4 72000_60000_M4 0.012
r 72000_60000_M4 76000_60000_M4 0.012
r 76000_60000_M4 80000_60000_M4 0.012
r 80000_60000_M4 84000_60000_M4 0.012
r 84000_60000_M4 88000_60000_M4 0.012
r 88000_60000_M4 92000_60000_M4 0.012
r 92000_60000_M4 96000_60000_M4 0.012
r 96000_60000_M4 100000_60000_M4 0.012
r 4000_64000_M4 8000_64000_M4 0.012
r 8000_64000_M4 12000_64000_M4 0.012
r 12000_64000_M4 16000_64000_M4 0.012
r 16000_64000_M4 20000_64000_M4 0.012
r 20000_64000_M4 24000_64000_M4 0.012
r 24000_64000_M4 28000_64000_M4 0.012
r 28000_64000_M4 32000_64000_M4 0.012
r 32000_64000_M4 36000_64000_M4 0.012
r 36000_64000_M4 40000_64000_M4 0.012
r 40000_64000_M4 44000_64000_M4 0.012
r 44000_64000_M4 48000_64000_M4 0.012
r 48000_64000_M4 52000_64000_M4 0.012
r 52000_64000_M4 56000_64000_M4 0.012
r 56000_64000_M4 60000_64000_M4 0.012
r 60000_64000_M4 64000_64000_M4 0.012
r 64000_64000_M4 68000_64000_M4 0.012
r 68000_64000_M4 72000_64000_M4 0.012
r 72000_64000_M4 76000_64000_M4 0.012
r 76000_64000_M4 80000_64000_M4 0.012
r 80000_64000_M4 84000_64000_M4 0.012
r 84000_64000_M4 88000_64000_M4 0.012
r 88000_64000_M4 92000_64000_M4 0.012
r 92000_64000_M4 96000_64000_M4 0.012
r 96000_64000_M4 100000_64000_M4 0.012
r 4000_68000_M4 8000_68000_M4 0.012
r 8000_68000_M4 12000_68000_M4 0.012
r 12000_68000_M4 16000_68000_M4 0.012
r 16000_68000_M4 20000_68000_M4 0.012
r 20000_68000_M4 24000_68000_M4 0.012
r 24000_68000_M4 28000_68000_M4 0.012
r 28000_68000_M4 32000_68000_M4 0.012
r 32000_68000_M4 36000_68000_M4 0.012
r 36000_68000_M4 40000_68000_M4 0.012
r 40000_68000_M4 44000_68000_M4 0.012
r 44000_68000_M4 48000_68000_M4 0.012
r 48000_68000_M4 52000_68000_M4 0.012
r 52000_68000_M4 56000_68000_M4 0.012
r 56000_68000_M4 60000_68000_M4 0.012
r 60000_68000_M4 64000_68000_M4 0.012
r 64000_68000_M4 68000_68000_M4 0.012
r 68000_68000_M4 72000_68000_M4 0.012
r 72000_68000_M4 76000_68000_M4 0.012
r 76000_68000_M4 80000_68000_M4 0.012
r 80000_68000_M4 84000_68000_M4 0.012
r 84000_68000_M4 88000_68000_M4 0.012
r 88000_68000_M4 92000_68000_M4 0.012
r 92000_68000_M4 96000_68000_M4 0.012
r 96000_68000_M4 100000_68000_M4 0.012
r 4000_72000_M4 8000_72000_M4 0.012
r 8000_72000_M4 12000_72000_M4 0.012
r 12000_72000_M4 16000_72000_M4 0.012
r 16000_72000_M4 20000_72000_M4 0.012
r 20000_72000_M4 24000_72000_M4 0.012
r 24000_72000_M4 28000_72000_M4 0.012
r 28000_72000_M4 32000_72000_M4 0.012
r 32000_72000_M4 36000_72000_M4 0.012
r 36000_72000_M4 40000_72000_M4 0.012
r 40000_72000_M4 44000_72000_M4 0.012
r 44000_72000_M4 48000_72000_M4 0.012
r 48000_72000_M4 52000_72000_M4 0.012
r 52000_72000_M4 56000_72000_M4 0.012
r 56000_72000_M4 60000_72000_M4 0.012
r 60000_72000_M4 64000_72000_M4 0.012
r 64000_72000_M4 68000_72000_M4 0.012
r 68000_72000_M4 72000_72000_M4 0.012
r 72000_72000_M4 76000_72000_M4 0.012
r 76000_72000_M4 80000_72000_M4 0.012
r 80000_72000_M4 84000_72000_M4 0.012
r 84000_72000_M4 88000_72000_M4 0.012
r 88000_72000_M4 92000_72000_M4 0.012
r 92000_72000_M4 96000_72000_M4 0.012
r 96000_72000_M4 100000_72000_M4 0.012
r 4000_76000_M4 8000_76000_M4 0.012
r 8000_76000_M4 12000_76000_M4 0.012
r 12000_76000_M4 16000_76000_M4 0.012
r 16000_76000_M4 20000_76000_M4 0.012
r 20000_76000_M4 24000_76000_M4 0.012
r 24000_76000_M4 28000_76000_M4 0.012
r 28000_76000_M4 32000_76000_M4 0.012
r 32000_76000_M4 36000_76000_M4 0.012
r 36000_76000_M4 40000_76000_M4 0.012
r 40000_76000_M4 44000_76000_M4 0.012
r 44000_76000_M4 48000_76000_M4 0.012
r 48000_76000_M4 52000_76000_M4 0.012
r 52000_76000_M4 56000_76000_M4 0.012
r 56000_76000_M4 60000_76000_M4 0.012
r 60000_76000_M4 64000_76000_M4 0.012
r 64000_76000_M4 68000_76000_M4 0.012
r 68000_76000_M4 72000_76000_M4 0.012
r 72000_76000_M4 76000_76000_M4 0.012
r 76000_76000_M4 80000_76000_M4 0.012
r 80000_76000_M4 84000_76000_M4 0.012
r 84000_76000_M4 88000_76000_M4 0.012
r 88000_76000_M4 92000_76000_M4 0.012
r 92000_76000_M4 96000_76000_M4 0.012
r 96000_76000_M4 100000_76000_M4 0.012
r 4000_80000_M4 8000_80000_M4 0.012
r 8000_80000_M4 12000_80000_M4 0.012
r 12000_80000_M4 16000_80000_M4 0.012
r 16000_80000_M4 20000_80000_M4 0.012
r 20000_80000_M4 24000_80000_M4 0.012
r 24000_80000_M4 28000_80000_M4 0.012
r 28000_80000_M4 32000_80000_M4 0.012
r 32000_80000_M4 36000_80000_M4 0.012
r 36000_80000_M4 40000_80000_M4 0.012
r 40000_80000_M4 44000_80000_M4 0.012
r 44000_80000_M4 48000_80000_M4 0.012
r 48000_80000_M4 52000_80000_M4 0.012
r 52000_80000_M4 56000_80000_M4 0.012
r 56000_80000_M4 60000_80000_M4 0.012
r 60000_80000_M4 64000_80000_M4 0.012
r 64000_80000_M4 68000_80000_M4 0.012
r 68000_80000_M4 72000_80000_M4 0.012
r 72000_80000_M4 76000_80000_M4 0.012
r 76000_80000_M4 80000_80000_M4 0.012
r 80000_80000_M4 84000_80000_M4 0.012
r 84000_80000_M4 88000_80000_M4 0.012
r 88000_80000_M4 92000_80000_M4 0.012
r 92000_80000_M4 96000_80000_M4 0.012
r 96000_80000_M4 100000_80000_M4 0.012
r 4000_84000_M4 8000_84000_M4 0.012
r 8000_84000_M4 12000_84000_M4 0.012
r 12000_84000_M4 16000_84000_M4 0.012
r 16000_84000_M4 20000_84000_M4 0.012
r 20000_84000_M4 24000_84000_M4 0.012
r 24000_84000_M4 28000_84000_M4 0.012
r 28000_84000_M4 32000_84000_M4 0.012
r 32000_84000_M4 36000_84000_M4 0.012
r 36000_84000_M4 40000_84000_M4 0.012
r 40000_84000_M4 44000_84000_M4 0.012
r 44000_84000_M4 48000_84000_M4 0.012
r 48000_84000_M4 52000_84000_M4 0.012
r 52000_84000_M4 56000_84000_M4 0.012
r 56000_84000_M4 60000_84000_M4 0.012
r 60000_84000_M4 64000_84000_M4 0.012
r 64000_84000_M4 68000_84000_M4 0.012
r 68000_84000_M4 72000_84000_M4 0.012
r 72000_84000_M4 76000_84000_M4 0.012
r 76000_84000_M4 80000_84000_M4 0.012
r 80000_84000_M4 84000_84000_M4 0.012
r 84000_84000_M4 88000_84000_M4 0.012
r 88000_84000_M4 92000_84000_M4 0.012
r 92000_84000_M4 96000_84000_M4 0.012
r 96000_84000_M4 100000_84000_M4 0.012
r 4000_88000_M4 8000_88000_M4 0.012
r 8000_88000_M4 12000_88000_M4 0.012
r 12000_88000_M4 16000_88000_M4 0.012
r 16000_88000_M4 20000_88000_M4 0.012
r 20000_88000_M4 24000_88000_M4 0.012
r 24000_88000_M4 28000_88000_M4 0.012
r 28000_88000_M4 32000_88000_M4 0.012
r 32000_88000_M4 36000_88000_M4 0.012
r 36000_88000_M4 40000_88000_M4 0.012
r 40000_88000_M4 44000_88000_M4 0.012
r 44000_88000_M4 48000_88000_M4 0.012
r 48000_88000_M4 52000_88000_M4 0.012
r 52000_88000_M4 56000_88000_M4 0.012
r 56000_88000_M4 60000_88000_M4 0.012
r 60000_88000_M4 64000_88000_M4 0.012
r 64000_88000_M4 68000_88000_M4 0.012
r 68000_88000_M4 72000_88000_M4 0.012
r 72000_88000_M4 76000_88000_M4 0.012
r 76000_88000_M4 80000_88000_M4 0.012
r 80000_88000_M4 84000_88000_M4 0.012
r 84000_88000_M4 88000_88000_M4 0.012
r 88000_88000_M4 92000_88000_M4 0.012
r 92000_88000_M4 96000_88000_M4 0.012
r 96000_88000_M4 100000_88000_M4 0.012
r 4000_92000_M4 8000_92000_M4 0.012
r 8000_92000_M4 12000_92000_M4 0.012
r 12000_92000_M4 16000_92000_M4 0.012
r 16000_92000_M4 20000_92000_M4 0.012
r 20000_92000_M4 24000_92000_M4 0.012
r 24000_92000_M4 28000_92000_M4 0.012
r 28000_92000_M4 32000_92000_M4 0.012
r 32000_92000_M4 36000_92000_M4 0.012
r 36000_92000_M4 40000_92000_M4 0.012
r 40000_92000_M4 44000_92000_M4 0.012
r 44000_92000_M4 48000_92000_M4 0.012
r 48000_92000_M4 52000_92000_M4 0.012
r 52000_92000_M4 56000_92000_M4 0.012
r 56000_92000_M4 60000_92000_M4 0.012
r 60000_92000_M4 64000_92000_M4 0.012
r 64000_92000_M4 68000_92000_M4 0.012
r 68000_92000_M4 72000_92000_M4 0.012
r 72000_92000_M4 76000_92000_M4 0.012
r 76000_92000_M4 80000_92000_M4 0.012
r 80000_92000_M4 84000_92000_M4 0.012
r 84000_92000_M4 88000_92000_M4 0.012
r 88000_92000_M4 92000_92000_M4 0.012
r 92000_92000_M4 96000_92000_M4 0.012
r 96000_92000_M4 100000_92000_M4 0.012
r 4000_96000_M4 8000_96000_M4 0.012
r 8000_96000_M4 12000_96000_M4 0.012
r 12000_96000_M4 16000_96000_M4 0.012
r 16000_96000_M4 20000_96000_M4 0.012
r 20000_96000_M4 24000_96000_M4 0.012
r 24000_96000_M4 28000_96000_M4 0.012
r 28000_96000_M4 32000_96000_M4 0.012
r 32000_96000_M4 36000_96000_M4 0.012
r 36000_96000_M4 40000_96000_M4 0.012
r 40000_96000_M4 44000_96000_M4 0.012
r 44000_96000_M4 48000_96000_M4 0.012
r 48000_96000_M4 52000_96000_M4 0.012
r 52000_96000_M4 56000_96000_M4 0.012
r 56000_96000_M4 60000_96000_M4 0.012
r 60000_96000_M4 64000_96000_M4 0.012
r 64000_96000_M4 68000_96000_M4 0.012
r 68000_96000_M4 72000_96000_M4 0.012
r 72000_96000_M4 76000_96000_M4 0.012
r 76000_96000_M4 80000_96000_M4 0.012
r 80000_96000_M4 84000_96000_M4 0.012
r 84000_96000_M4 88000_96000_M4 0.012
r 88000_96000_M4 92000_96000_M4 0.012
r 92000_96000_M4 96000_96000_M4 0.012
r 96000_96000_M4 100000_96000_M4 0.012
r 4000_100000_M4 8000_100000_M4 0.012
r 8000_100000_M4 12000_100000_M4 0.012
r 12000_100000_M4 16000_100000_M4 0.012
r 16000_100000_M4 20000_100000_M4 0.012
r 20000_100000_M4 24000_100000_M4 0.012
r 24000_100000_M4 28000_100000_M4 0.012
r 28000_100000_M4 32000_100000_M4 0.012
r 32000_100000_M4 36000_100000_M4 0.012
r 36000_100000_M4 40000_100000_M4 0.012
r 40000_100000_M4 44000_100000_M4 0.012
r 44000_100000_M4 48000_100000_M4 0.012
r 48000_100000_M4 52000_100000_M4 0.012
r 52000_100000_M4 56000_100000_M4 0.012
r 56000_100000_M4 60000_100000_M4 0.012
r 60000_100000_M4 64000_100000_M4 0.012
r 64000_100000_M4 68000_100000_M4 0.012
r 68000_100000_M4 72000_100000_M4 0.012
r 72000_100000_M4 76000_100000_M4 0.012
r 76000_100000_M4 80000_100000_M4 0.012
r 80000_100000_M4 84000_100000_M4 0.012
r 84000_100000_M4 88000_100000_M4 0.012
r 88000_100000_M4 92000_100000_M4 0.012
r 92000_100000_M4 96000_100000_M4 0.012
r 96000_100000_M4 100000_100000_M4 0.012

* M4 Vertical resistors
r 4000_4000_M4 4000_8000_M4 0.015
r 4000_8000_M4 4000_12000_M4 0.015
r 4000_12000_M4 4000_16000_M4 0.015
r 4000_16000_M4 4000_20000_M4 0.015
r 4000_20000_M4 4000_24000_M4 0.015
r 4000_24000_M4 4000_28000_M4 0.015
r 4000_28000_M4 4000_32000_M4 0.015
r 4000_32000_M4 4000_36000_M4 0.015
r 4000_36000_M4 4000_40000_M4 0.015
r 4000_40000_M4 4000_44000_M4 0.015
r 4000_44000_M4 4000_48000_M4 0.015
r 4000_48000_M4 4000_52000_M4 0.015
r 4000_52000_M4 4000_56000_M4 0.015
r 4000_56000_M4 4000_60000_M4 0.015
r 4000_60000_M4 4000_64000_M4 0.015
r 4000_64000_M4 4000_68000_M4 0.015
r 4000_68000_M4 4000_72000_M4 0.015
r 4000_72000_M4 4000_76000_M4 0.015
r 4000_76000_M4 4000_80000_M4 0.015
r 4000_80000_M4 4000_84000_M4 0.015
r 4000_84000_M4 4000_88000_M4 0.015
r 4000_88000_M4 4000_92000_M4 0.015
r 4000_92000_M4 4000_96000_M4 0.015
r 4000_96000_M4 4000_100000_M4 0.015
r 8000_4000_M4 8000_8000_M4 0.015
r 8000_8000_M4 8000_12000_M4 0.015
r 8000_12000_M4 8000_16000_M4 0.015
r 8000_16000_M4 8000_20000_M4 0.015
r 8000_20000_M4 8000_24000_M4 0.015
r 8000_24000_M4 8000_28000_M4 0.015
r 8000_28000_M4 8000_32000_M4 0.015
r 8000_32000_M4 8000_36000_M4 0.015
r 8000_36000_M4 8000_40000_M4 0.015
r 8000_40000_M4 8000_44000_M4 0.015
r 8000_44000_M4 8000_48000_M4 0.015
r 8000_48000_M4 8000_52000_M4 0.015
r 8000_52000_M4 8000_56000_M4 0.015
r 8000_56000_M4 8000_60000_M4 0.015
r 8000_60000_M4 8000_64000_M4 0.015
r 8000_64000_M4 8000_68000_M4 0.015
r 8000_68000_M4 8000_72000_M4 0.015
r 8000_72000_M4 8000_76000_M4 0.015
r 8000_76000_M4 8000_80000_M4 0.015
r 8000_80000_M4 8000_84000_M4 0.015
r 8000_84000_M4 8000_88000_M4 0.015
r 8000_88000_M4 8000_92000_M4 0.015
r 8000_92000_M4 8000_96000_M4 0.015
r 8000_96000_M4 8000_100000_M4 0.015
r 12000_4000_M4 12000_8000_M4 0.015
r 12000_8000_M4 12000_12000_M4 0.015
r 12000_12000_M4 12000_16000_M4 0.015
r 12000_16000_M4 12000_20000_M4 0.015
r 12000_20000_M4 12000_24000_M4 0.015
r 12000_24000_M4 12000_28000_M4 0.015
r 12000_28000_M4 12000_32000_M4 0.015
r 12000_32000_M4 12000_36000_M4 0.015
r 12000_36000_M4 12000_40000_M4 0.015
r 12000_40000_M4 12000_44000_M4 0.015
r 12000_44000_M4 12000_48000_M4 0.015
r 12000_48000_M4 12000_52000_M4 0.015
r 12000_52000_M4 12000_56000_M4 0.015
r 12000_56000_M4 12000_60000_M4 0.015
r 12000_60000_M4 12000_64000_M4 0.015
r 12000_64000_M4 12000_68000_M4 0.015
r 12000_68000_M4 12000_72000_M4 0.015
r 12000_72000_M4 12000_76000_M4 0.015
r 12000_76000_M4 12000_80000_M4 0.015
r 12000_80000_M4 12000_84000_M4 0.015
r 12000_84000_M4 12000_88000_M4 0.015
r 12000_88000_M4 12000_92000_M4 0.015
r 12000_92000_M4 12000_96000_M4 0.015
r 12000_96000_M4 12000_100000_M4 0.015
r 16000_4000_M4 16000_8000_M4 0.015
r 16000_8000_M4 16000_12000_M4 0.015
r 16000_12000_M4 16000_16000_M4 0.015
r 16000_16000_M4 16000_20000_M4 0.015
r 16000_20000_M4 16000_24000_M4 0.015
r 16000_24000_M4 16000_28000_M4 0.015
r 16000_28000_M4 16000_32000_M4 0.015
r 16000_32000_M4 16000_36000_M4 0.015
r 16000_36000_M4 16000_40000_M4 0.015
r 16000_40000_M4 16000_44000_M4 0.015
r 16000_44000_M4 16000_48000_M4 0.015
r 16000_48000_M4 16000_52000_M4 0.015
r 16000_52000_M4 16000_56000_M4 0.015
r 16000_56000_M4 16000_60000_M4 0.015
r 16000_60000_M4 16000_64000_M4 0.015
r 16000_64000_M4 16000_68000_M4 0.015
r 16000_68000_M4 16000_72000_M4 0.015
r 16000_72000_M4 16000_76000_M4 0.015
r 16000_76000_M4 16000_80000_M4 0.015
r 16000_80000_M4 16000_84000_M4 0.015
r 16000_84000_M4 16000_88000_M4 0.015
r 16000_88000_M4 16000_92000_M4 0.015
r 16000_92000_M4 16000_96000_M4 0.015
r 16000_96000_M4 16000_100000_M4 0.015
r 20000_4000_M4 20000_8000_M4 0.015
r 20000_8000_M4 20000_12000_M4 0.015
r 20000_12000_M4 20000_16000_M4 0.015
r 20000_16000_M4 20000_20000_M4 0.015
r 20000_20000_M4 20000_24000_M4 0.015
r 20000_24000_M4 20000_28000_M4 0.015
r 20000_28000_M4 20000_32000_M4 0.015
r 20000_32000_M4 20000_36000_M4 0.015
r 20000_36000_M4 20000_40000_M4 0.015
r 20000_40000_M4 20000_44000_M4 0.015
r 20000_44000_M4 20000_48000_M4 0.015
r 20000_48000_M4 20000_52000_M4 0.015
r 20000_52000_M4 20000_56000_M4 0.015
r 20000_56000_M4 20000_60000_M4 0.015
r 20000_60000_M4 20000_64000_M4 0.015
r 20000_64000_M4 20000_68000_M4 0.015
r 20000_68000_M4 20000_72000_M4 0.015
r 20000_72000_M4 20000_76000_M4 0.015
r 20000_76000_M4 20000_80000_M4 0.015
r 20000_80000_M4 20000_84000_M4 0.015
r 20000_84000_M4 20000_88000_M4 0.015
r 20000_88000_M4 20000_92000_M4 0.015
r 20000_92000_M4 20000_96000_M4 0.015
r 20000_96000_M4 20000_100000_M4 0.015
r 24000_4000_M4 24000_8000_M4 0.015
r 24000_8000_M4 24000_12000_M4 0.015
r 24000_12000_M4 24000_16000_M4 0.015
r 24000_16000_M4 24000_20000_M4 0.015
r 24000_20000_M4 24000_24000_M4 0.015
r 24000_24000_M4 24000_28000_M4 0.015
r 24000_28000_M4 24000_32000_M4 0.015
r 24000_32000_M4 24000_36000_M4 0.015
r 24000_36000_M4 24000_40000_M4 0.015
r 24000_40000_M4 24000_44000_M4 0.015
r 24000_44000_M4 24000_48000_M4 0.015
r 24000_48000_M4 24000_52000_M4 0.015
r 24000_52000_M4 24000_56000_M4 0.015
r 24000_56000_M4 24000_60000_M4 0.015
r 24000_60000_M4 24000_64000_M4 0.015
r 24000_64000_M4 24000_68000_M4 0.015
r 24000_68000_M4 24000_72000_M4 0.015
r 24000_72000_M4 24000_76000_M4 0.015
r 24000_76000_M4 24000_80000_M4 0.015
r 24000_80000_M4 24000_84000_M4 0.015
r 24000_84000_M4 24000_88000_M4 0.015
r 24000_88000_M4 24000_92000_M4 0.015
r 24000_92000_M4 24000_96000_M4 0.015
r 24000_96000_M4 24000_100000_M4 0.015
r 28000_4000_M4 28000_8000_M4 0.015
r 28000_8000_M4 28000_12000_M4 0.015
r 28000_12000_M4 28000_16000_M4 0.015
r 28000_16000_M4 28000_20000_M4 0.015
r 28000_20000_M4 28000_24000_M4 0.015
r 28000_24000_M4 28000_28000_M4 0.015
r 28000_28000_M4 28000_32000_M4 0.015
r 28000_32000_M4 28000_36000_M4 0.015
r 28000_36000_M4 28000_40000_M4 0.015
r 28000_40000_M4 28000_44000_M4 0.015
r 28000_44000_M4 28000_48000_M4 0.015
r 28000_48000_M4 28000_52000_M4 0.015
r 28000_52000_M4 28000_56000_M4 0.015
r 28000_56000_M4 28000_60000_M4 0.015
r 28000_60000_M4 28000_64000_M4 0.015
r 28000_64000_M4 28000_68000_M4 0.015
r 28000_68000_M4 28000_72000_M4 0.015
r 28000_72000_M4 28000_76000_M4 0.015
r 28000_76000_M4 28000_80000_M4 0.015
r 28000_80000_M4 28000_84000_M4 0.015
r 28000_84000_M4 28000_88000_M4 0.015
r 28000_88000_M4 28000_92000_M4 0.015
r 28000_92000_M4 28000_96000_M4 0.015
r 28000_96000_M4 28000_100000_M4 0.015
r 32000_4000_M4 32000_8000_M4 0.015
r 32000_8000_M4 32000_12000_M4 0.015
r 32000_12000_M4 32000_16000_M4 0.015
r 32000_16000_M4 32000_20000_M4 0.015
r 32000_20000_M4 32000_24000_M4 0.015
r 32000_24000_M4 32000_28000_M4 0.015
r 32000_28000_M4 32000_32000_M4 0.015
r 32000_32000_M4 32000_36000_M4 0.015
r 32000_36000_M4 32000_40000_M4 0.015
r 32000_40000_M4 32000_44000_M4 0.015
r 32000_44000_M4 32000_48000_M4 0.015
r 32000_48000_M4 32000_52000_M4 0.015
r 32000_52000_M4 32000_56000_M4 0.015
r 32000_56000_M4 32000_60000_M4 0.015
r 32000_60000_M4 32000_64000_M4 0.015
r 32000_64000_M4 32000_68000_M4 0.015
r 32000_68000_M4 32000_72000_M4 0.015
r 32000_72000_M4 32000_76000_M4 0.015
r 32000_76000_M4 32000_80000_M4 0.015
r 32000_80000_M4 32000_84000_M4 0.015
r 32000_84000_M4 32000_88000_M4 0.015
r 32000_88000_M4 32000_92000_M4 0.015
r 32000_92000_M4 32000_96000_M4 0.015
r 32000_96000_M4 32000_100000_M4 0.015
r 36000_4000_M4 36000_8000_M4 0.015
r 36000_8000_M4 36000_12000_M4 0.015
r 36000_12000_M4 36000_16000_M4 0.015
r 36000_16000_M4 36000_20000_M4 0.015
r 36000_20000_M4 36000_24000_M4 0.015
r 36000_24000_M4 36000_28000_M4 0.015
r 36000_28000_M4 36000_32000_M4 0.015
r 36000_32000_M4 36000_36000_M4 0.015
r 36000_36000_M4 36000_40000_M4 0.015
r 36000_40000_M4 36000_44000_M4 0.015
r 36000_44000_M4 36000_48000_M4 0.015
r 36000_48000_M4 36000_52000_M4 0.015
r 36000_52000_M4 36000_56000_M4 0.015
r 36000_56000_M4 36000_60000_M4 0.015
r 36000_60000_M4 36000_64000_M4 0.015
r 36000_64000_M4 36000_68000_M4 0.015
r 36000_68000_M4 36000_72000_M4 0.015
r 36000_72000_M4 36000_76000_M4 0.015
r 36000_76000_M4 36000_80000_M4 0.015
r 36000_80000_M4 36000_84000_M4 0.015
r 36000_84000_M4 36000_88000_M4 0.015
r 36000_88000_M4 36000_92000_M4 0.015
r 36000_92000_M4 36000_96000_M4 0.015
r 36000_96000_M4 36000_100000_M4 0.015
r 40000_4000_M4 40000_8000_M4 0.015
r 40000_8000_M4 40000_12000_M4 0.015
r 40000_12000_M4 40000_16000_M4 0.015
r 40000_16000_M4 40000_20000_M4 0.015
r 40000_20000_M4 40000_24000_M4 0.015
r 40000_24000_M4 40000_28000_M4 0.015
r 40000_28000_M4 40000_32000_M4 0.015
r 40000_32000_M4 40000_36000_M4 0.015
r 40000_36000_M4 40000_40000_M4 0.015
r 40000_40000_M4 40000_44000_M4 0.015
r 40000_44000_M4 40000_48000_M4 0.015
r 40000_48000_M4 40000_52000_M4 0.015
r 40000_52000_M4 40000_56000_M4 0.015
r 40000_56000_M4 40000_60000_M4 0.015
r 40000_60000_M4 40000_64000_M4 0.015
r 40000_64000_M4 40000_68000_M4 0.015
r 40000_68000_M4 40000_72000_M4 0.015
r 40000_72000_M4 40000_76000_M4 0.015
r 40000_76000_M4 40000_80000_M4 0.015
r 40000_80000_M4 40000_84000_M4 0.015
r 40000_84000_M4 40000_88000_M4 0.015
r 40000_88000_M4 40000_92000_M4 0.015
r 40000_92000_M4 40000_96000_M4 0.015
r 40000_96000_M4 40000_100000_M4 0.015
r 44000_4000_M4 44000_8000_M4 0.015
r 44000_8000_M4 44000_12000_M4 0.015
r 44000_12000_M4 44000_16000_M4 0.015
r 44000_16000_M4 44000_20000_M4 0.015
r 44000_20000_M4 44000_24000_M4 0.015
r 44000_24000_M4 44000_28000_M4 0.015
r 44000_28000_M4 44000_32000_M4 0.015
r 44000_32000_M4 44000_36000_M4 0.015
r 44000_36000_M4 44000_40000_M4 0.015
r 44000_40000_M4 44000_44000_M4 0.015
r 44000_44000_M4 44000_48000_M4 0.015
r 44000_48000_M4 44000_52000_M4 0.015
r 44000_52000_M4 44000_56000_M4 0.015
r 44000_56000_M4 44000_60000_M4 0.015
r 44000_60000_M4 44000_64000_M4 0.015
r 44000_64000_M4 44000_68000_M4 0.015
r 44000_68000_M4 44000_72000_M4 0.015
r 44000_72000_M4 44000_76000_M4 0.015
r 44000_76000_M4 44000_80000_M4 0.015
r 44000_80000_M4 44000_84000_M4 0.015
r 44000_84000_M4 44000_88000_M4 0.015
r 44000_88000_M4 44000_92000_M4 0.015
r 44000_92000_M4 44000_96000_M4 0.015
r 44000_96000_M4 44000_100000_M4 0.015
r 48000_4000_M4 48000_8000_M4 0.015
r 48000_8000_M4 48000_12000_M4 0.015
r 48000_12000_M4 48000_16000_M4 0.015
r 48000_16000_M4 48000_20000_M4 0.015
r 48000_20000_M4 48000_24000_M4 0.015
r 48000_24000_M4 48000_28000_M4 0.015
r 48000_28000_M4 48000_32000_M4 0.015
r 48000_32000_M4 48000_36000_M4 0.015
r 48000_36000_M4 48000_40000_M4 0.015
r 48000_40000_M4 48000_44000_M4 0.015
r 48000_44000_M4 48000_48000_M4 0.015
r 48000_48000_M4 48000_52000_M4 0.015
r 48000_52000_M4 48000_56000_M4 0.015
r 48000_56000_M4 48000_60000_M4 0.015
r 48000_60000_M4 48000_64000_M4 0.015
r 48000_64000_M4 48000_68000_M4 0.015
r 48000_68000_M4 48000_72000_M4 0.015
r 48000_72000_M4 48000_76000_M4 0.015
r 48000_76000_M4 48000_80000_M4 0.015
r 48000_80000_M4 48000_84000_M4 0.015
r 48000_84000_M4 48000_88000_M4 0.015
r 48000_88000_M4 48000_92000_M4 0.015
r 48000_92000_M4 48000_96000_M4 0.015
r 48000_96000_M4 48000_100000_M4 0.015
r 52000_4000_M4 52000_8000_M4 0.015
r 52000_8000_M4 52000_12000_M4 0.015
r 52000_12000_M4 52000_16000_M4 0.015
r 52000_16000_M4 52000_20000_M4 0.015
r 52000_20000_M4 52000_24000_M4 0.015
r 52000_24000_M4 52000_28000_M4 0.015
r 52000_28000_M4 52000_32000_M4 0.015
r 52000_32000_M4 52000_36000_M4 0.015
r 52000_36000_M4 52000_40000_M4 0.015
r 52000_40000_M4 52000_44000_M4 0.015
r 52000_44000_M4 52000_48000_M4 0.015
r 52000_48000_M4 52000_52000_M4 0.015
r 52000_52000_M4 52000_56000_M4 0.015
r 52000_56000_M4 52000_60000_M4 0.015
r 52000_60000_M4 52000_64000_M4 0.015
r 52000_64000_M4 52000_68000_M4 0.015
r 52000_68000_M4 52000_72000_M4 0.015
r 52000_72000_M4 52000_76000_M4 0.015
r 52000_76000_M4 52000_80000_M4 0.015
r 52000_80000_M4 52000_84000_M4 0.015
r 52000_84000_M4 52000_88000_M4 0.015
r 52000_88000_M4 52000_92000_M4 0.015
r 52000_92000_M4 52000_96000_M4 0.015
r 52000_96000_M4 52000_100000_M4 0.015
r 56000_4000_M4 56000_8000_M4 0.015
r 56000_8000_M4 56000_12000_M4 0.015
r 56000_12000_M4 56000_16000_M4 0.015
r 56000_16000_M4 56000_20000_M4 0.015
r 56000_20000_M4 56000_24000_M4 0.015
r 56000_24000_M4 56000_28000_M4 0.015
r 56000_28000_M4 56000_32000_M4 0.015
r 56000_32000_M4 56000_36000_M4 0.015
r 56000_36000_M4 56000_40000_M4 0.015
r 56000_40000_M4 56000_44000_M4 0.015
r 56000_44000_M4 56000_48000_M4 0.015
r 56000_48000_M4 56000_52000_M4 0.015
r 56000_52000_M4 56000_56000_M4 0.015
r 56000_56000_M4 56000_60000_M4 0.015
r 56000_60000_M4 56000_64000_M4 0.015
r 56000_64000_M4 56000_68000_M4 0.015
r 56000_68000_M4 56000_72000_M4 0.015
r 56000_72000_M4 56000_76000_M4 0.015
r 56000_76000_M4 56000_80000_M4 0.015
r 56000_80000_M4 56000_84000_M4 0.015
r 56000_84000_M4 56000_88000_M4 0.015
r 56000_88000_M4 56000_92000_M4 0.015
r 56000_92000_M4 56000_96000_M4 0.015
r 56000_96000_M4 56000_100000_M4 0.015
r 60000_4000_M4 60000_8000_M4 0.015
r 60000_8000_M4 60000_12000_M4 0.015
r 60000_12000_M4 60000_16000_M4 0.015
r 60000_16000_M4 60000_20000_M4 0.015
r 60000_20000_M4 60000_24000_M4 0.015
r 60000_24000_M4 60000_28000_M4 0.015
r 60000_28000_M4 60000_32000_M4 0.015
r 60000_32000_M4 60000_36000_M4 0.015
r 60000_36000_M4 60000_40000_M4 0.015
r 60000_40000_M4 60000_44000_M4 0.015
r 60000_44000_M4 60000_48000_M4 0.015
r 60000_48000_M4 60000_52000_M4 0.015
r 60000_52000_M4 60000_56000_M4 0.015
r 60000_56000_M4 60000_60000_M4 0.015
r 60000_60000_M4 60000_64000_M4 0.015
r 60000_64000_M4 60000_68000_M4 0.015
r 60000_68000_M4 60000_72000_M4 0.015
r 60000_72000_M4 60000_76000_M4 0.015
r 60000_76000_M4 60000_80000_M4 0.015
r 60000_80000_M4 60000_84000_M4 0.015
r 60000_84000_M4 60000_88000_M4 0.015
r 60000_88000_M4 60000_92000_M4 0.015
r 60000_92000_M4 60000_96000_M4 0.015
r 60000_96000_M4 60000_100000_M4 0.015
r 64000_4000_M4 64000_8000_M4 0.015
r 64000_8000_M4 64000_12000_M4 0.015
r 64000_12000_M4 64000_16000_M4 0.015
r 64000_16000_M4 64000_20000_M4 0.015
r 64000_20000_M4 64000_24000_M4 0.015
r 64000_24000_M4 64000_28000_M4 0.015
r 64000_28000_M4 64000_32000_M4 0.015
r 64000_32000_M4 64000_36000_M4 0.015
r 64000_36000_M4 64000_40000_M4 0.015
r 64000_40000_M4 64000_44000_M4 0.015
r 64000_44000_M4 64000_48000_M4 0.015
r 64000_48000_M4 64000_52000_M4 0.015
r 64000_52000_M4 64000_56000_M4 0.015
r 64000_56000_M4 64000_60000_M4 0.015
r 64000_60000_M4 64000_64000_M4 0.015
r 64000_64000_M4 64000_68000_M4 0.015
r 64000_68000_M4 64000_72000_M4 0.015
r 64000_72000_M4 64000_76000_M4 0.015
r 64000_76000_M4 64000_80000_M4 0.015
r 64000_80000_M4 64000_84000_M4 0.015
r 64000_84000_M4 64000_88000_M4 0.015
r 64000_88000_M4 64000_92000_M4 0.015
r 64000_92000_M4 64000_96000_M4 0.015
r 64000_96000_M4 64000_100000_M4 0.015
r 68000_4000_M4 68000_8000_M4 0.015
r 68000_8000_M4 68000_12000_M4 0.015
r 68000_12000_M4 68000_16000_M4 0.015
r 68000_16000_M4 68000_20000_M4 0.015
r 68000_20000_M4 68000_24000_M4 0.015
r 68000_24000_M4 68000_28000_M4 0.015
r 68000_28000_M4 68000_32000_M4 0.015
r 68000_32000_M4 68000_36000_M4 0.015
r 68000_36000_M4 68000_40000_M4 0.015
r 68000_40000_M4 68000_44000_M4 0.015
r 68000_44000_M4 68000_48000_M4 0.015
r 68000_48000_M4 68000_52000_M4 0.015
r 68000_52000_M4 68000_56000_M4 0.015
r 68000_56000_M4 68000_60000_M4 0.015
r 68000_60000_M4 68000_64000_M4 0.015
r 68000_64000_M4 68000_68000_M4 0.015
r 68000_68000_M4 68000_72000_M4 0.015
r 68000_72000_M4 68000_76000_M4 0.015
r 68000_76000_M4 68000_80000_M4 0.015
r 68000_80000_M4 68000_84000_M4 0.015
r 68000_84000_M4 68000_88000_M4 0.015
r 68000_88000_M4 68000_92000_M4 0.015
r 68000_92000_M4 68000_96000_M4 0.015
r 68000_96000_M4 68000_100000_M4 0.015
r 72000_4000_M4 72000_8000_M4 0.015
r 72000_8000_M4 72000_12000_M4 0.015
r 72000_12000_M4 72000_16000_M4 0.015
r 72000_16000_M4 72000_20000_M4 0.015
r 72000_20000_M4 72000_24000_M4 0.015
r 72000_24000_M4 72000_28000_M4 0.015
r 72000_28000_M4 72000_32000_M4 0.015
r 72000_32000_M4 72000_36000_M4 0.015
r 72000_36000_M4 72000_40000_M4 0.015
r 72000_40000_M4 72000_44000_M4 0.015
r 72000_44000_M4 72000_48000_M4 0.015
r 72000_48000_M4 72000_52000_M4 0.015
r 72000_52000_M4 72000_56000_M4 0.015
r 72000_56000_M4 72000_60000_M4 0.015
r 72000_60000_M4 72000_64000_M4 0.015
r 72000_64000_M4 72000_68000_M4 0.015
r 72000_68000_M4 72000_72000_M4 0.015
r 72000_72000_M4 72000_76000_M4 0.015
r 72000_76000_M4 72000_80000_M4 0.015
r 72000_80000_M4 72000_84000_M4 0.015
r 72000_84000_M4 72000_88000_M4 0.015
r 72000_88000_M4 72000_92000_M4 0.015
r 72000_92000_M4 72000_96000_M4 0.015
r 72000_96000_M4 72000_100000_M4 0.015
r 76000_4000_M4 76000_8000_M4 0.015
r 76000_8000_M4 76000_12000_M4 0.015
r 76000_12000_M4 76000_16000_M4 0.015
r 76000_16000_M4 76000_20000_M4 0.015
r 76000_20000_M4 76000_24000_M4 0.015
r 76000_24000_M4 76000_28000_M4 0.015
r 76000_28000_M4 76000_32000_M4 0.015
r 76000_32000_M4 76000_36000_M4 0.015
r 76000_36000_M4 76000_40000_M4 0.015
r 76000_40000_M4 76000_44000_M4 0.015
r 76000_44000_M4 76000_48000_M4 0.015
r 76000_48000_M4 76000_52000_M4 0.015
r 76000_52000_M4 76000_56000_M4 0.015
r 76000_56000_M4 76000_60000_M4 0.015
r 76000_60000_M4 76000_64000_M4 0.015
r 76000_64000_M4 76000_68000_M4 0.015
r 76000_68000_M4 76000_72000_M4 0.015
r 76000_72000_M4 76000_76000_M4 0.015
r 76000_76000_M4 76000_80000_M4 0.015
r 76000_80000_M4 76000_84000_M4 0.015
r 76000_84000_M4 76000_88000_M4 0.015
r 76000_88000_M4 76000_92000_M4 0.015
r 76000_92000_M4 76000_96000_M4 0.015
r 76000_96000_M4 76000_100000_M4 0.015
r 80000_4000_M4 80000_8000_M4 0.015
r 80000_8000_M4 80000_12000_M4 0.015
r 80000_12000_M4 80000_16000_M4 0.015
r 80000_16000_M4 80000_20000_M4 0.015
r 80000_20000_M4 80000_24000_M4 0.015
r 80000_24000_M4 80000_28000_M4 0.015
r 80000_28000_M4 80000_32000_M4 0.015
r 80000_32000_M4 80000_36000_M4 0.015
r 80000_36000_M4 80000_40000_M4 0.015
r 80000_40000_M4 80000_44000_M4 0.015
r 80000_44000_M4 80000_48000_M4 0.015
r 80000_48000_M4 80000_52000_M4 0.015
r 80000_52000_M4 80000_56000_M4 0.015
r 80000_56000_M4 80000_60000_M4 0.015
r 80000_60000_M4 80000_64000_M4 0.015
r 80000_64000_M4 80000_68000_M4 0.015
r 80000_68000_M4 80000_72000_M4 0.015
r 80000_72000_M4 80000_76000_M4 0.015
r 80000_76000_M4 80000_80000_M4 0.015
r 80000_80000_M4 80000_84000_M4 0.015
r 80000_84000_M4 80000_88000_M4 0.015
r 80000_88000_M4 80000_92000_M4 0.015
r 80000_92000_M4 80000_96000_M4 0.015
r 80000_96000_M4 80000_100000_M4 0.015
r 84000_4000_M4 84000_8000_M4 0.015
r 84000_8000_M4 84000_12000_M4 0.015
r 84000_12000_M4 84000_16000_M4 0.015
r 84000_16000_M4 84000_20000_M4 0.015
r 84000_20000_M4 84000_24000_M4 0.015
r 84000_24000_M4 84000_28000_M4 0.015
r 84000_28000_M4 84000_32000_M4 0.015
r 84000_32000_M4 84000_36000_M4 0.015
r 84000_36000_M4 84000_40000_M4 0.015
r 84000_40000_M4 84000_44000_M4 0.015
r 84000_44000_M4 84000_48000_M4 0.015
r 84000_48000_M4 84000_52000_M4 0.015
r 84000_52000_M4 84000_56000_M4 0.015
r 84000_56000_M4 84000_60000_M4 0.015
r 84000_60000_M4 84000_64000_M4 0.015
r 84000_64000_M4 84000_68000_M4 0.015
r 84000_68000_M4 84000_72000_M4 0.015
r 84000_72000_M4 84000_76000_M4 0.015
r 84000_76000_M4 84000_80000_M4 0.015
r 84000_80000_M4 84000_84000_M4 0.015
r 84000_84000_M4 84000_88000_M4 0.015
r 84000_88000_M4 84000_92000_M4 0.015
r 84000_92000_M4 84000_96000_M4 0.015
r 84000_96000_M4 84000_100000_M4 0.015
r 88000_4000_M4 88000_8000_M4 0.015
r 88000_8000_M4 88000_12000_M4 0.015
r 88000_12000_M4 88000_16000_M4 0.015
r 88000_16000_M4 88000_20000_M4 0.015
r 88000_20000_M4 88000_24000_M4 0.015
r 88000_24000_M4 88000_28000_M4 0.015
r 88000_28000_M4 88000_32000_M4 0.015
r 88000_32000_M4 88000_36000_M4 0.015
r 88000_36000_M4 88000_40000_M4 0.015
r 88000_40000_M4 88000_44000_M4 0.015
r 88000_44000_M4 88000_48000_M4 0.015
r 88000_48000_M4 88000_52000_M4 0.015
r 88000_52000_M4 88000_56000_M4 0.015
r 88000_56000_M4 88000_60000_M4 0.015
r 88000_60000_M4 88000_64000_M4 0.015
r 88000_64000_M4 88000_68000_M4 0.015
r 88000_68000_M4 88000_72000_M4 0.015
r 88000_72000_M4 88000_76000_M4 0.015
r 88000_76000_M4 88000_80000_M4 0.015
r 88000_80000_M4 88000_84000_M4 0.015
r 88000_84000_M4 88000_88000_M4 0.015
r 88000_88000_M4 88000_92000_M4 0.015
r 88000_92000_M4 88000_96000_M4 0.015
r 88000_96000_M4 88000_100000_M4 0.015
r 92000_4000_M4 92000_8000_M4 0.015
r 92000_8000_M4 92000_12000_M4 0.015
r 92000_12000_M4 92000_16000_M4 0.015
r 92000_16000_M4 92000_20000_M4 0.015
r 92000_20000_M4 92000_24000_M4 0.015
r 92000_24000_M4 92000_28000_M4 0.015
r 92000_28000_M4 92000_32000_M4 0.015
r 92000_32000_M4 92000_36000_M4 0.015
r 92000_36000_M4 92000_40000_M4 0.015
r 92000_40000_M4 92000_44000_M4 0.015
r 92000_44000_M4 92000_48000_M4 0.015
r 92000_48000_M4 92000_52000_M4 0.015
r 92000_52000_M4 92000_56000_M4 0.015
r 92000_56000_M4 92000_60000_M4 0.015
r 92000_60000_M4 92000_64000_M4 0.015
r 92000_64000_M4 92000_68000_M4 0.015
r 92000_68000_M4 92000_72000_M4 0.015
r 92000_72000_M4 92000_76000_M4 0.015
r 92000_76000_M4 92000_80000_M4 0.015
r 92000_80000_M4 92000_84000_M4 0.015
r 92000_84000_M4 92000_88000_M4 0.015
r 92000_88000_M4 92000_92000_M4 0.015
r 92000_92000_M4 92000_96000_M4 0.015
r 92000_96000_M4 92000_100000_M4 0.015
r 96000_4000_M4 96000_8000_M4 0.015
r 96000_8000_M4 96000_12000_M4 0.015
r 96000_12000_M4 96000_16000_M4 0.015
r 96000_16000_M4 96000_20000_M4 0.015
r 96000_20000_M4 96000_24000_M4 0.015
r 96000_24000_M4 96000_28000_M4 0.015
r 96000_28000_M4 96000_32000_M4 0.015
r 96000_32000_M4 96000_36000_M4 0.015
r 96000_36000_M4 96000_40000_M4 0.015
r 96000_40000_M4 96000_44000_M4 0.015
r 96000_44000_M4 96000_48000_M4 0.015
r 96000_48000_M4 96000_52000_M4 0.015
r 96000_52000_M4 96000_56000_M4 0.015
r 96000_56000_M4 96000_60000_M4 0.015
r 96000_60000_M4 96000_64000_M4 0.015
r 96000_64000_M4 96000_68000_M4 0.015
r 96000_68000_M4 96000_72000_M4 0.015
r 96000_72000_M4 96000_76000_M4 0.015
r 96000_76000_M4 96000_80000_M4 0.015
r 96000_80000_M4 96000_84000_M4 0.015
r 96000_84000_M4 96000_88000_M4 0.015
r 96000_88000_M4 96000_92000_M4 0.015
r 96000_92000_M4 96000_96000_M4 0.015
r 96000_96000_M4 96000_100000_M4 0.015
r 100000_4000_M4 100000_8000_M4 0.015
r 100000_8000_M4 100000_12000_M4 0.015
r 100000_12000_M4 100000_16000_M4 0.015
r 100000_16000_M4 100000_20000_M4 0.015
r 100000_20000_M4 100000_24000_M4 0.015
r 100000_24000_M4 100000_28000_M4 0.015
r 100000_28000_M4 100000_32000_M4 0.015
r 100000_32000_M4 100000_36000_M4 0.015
r 100000_36000_M4 100000_40000_M4 0.015
r 100000_40000_M4 100000_44000_M4 0.015
r 100000_44000_M4 100000_48000_M4 0.015
r 100000_48000_M4 100000_52000_M4 0.015
r 100000_52000_M4 100000_56000_M4 0.015
r 100000_56000_M4 100000_60000_M4 0.015
r 100000_60000_M4 100000_64000_M4 0.015
r 100000_64000_M4 100000_68000_M4 0.015
r 100000_68000_M4 100000_72000_M4 0.015
r 100000_72000_M4 100000_76000_M4 0.015
r 100000_76000_M4 100000_80000_M4 0.015
r 100000_80000_M4 100000_84000_M4 0.015
r 100000_84000_M4 100000_88000_M4 0.015
r 100000_88000_M4 100000_92000_M4 0.015
r 100000_92000_M4 100000_96000_M4 0.015
r 100000_96000_M4 100000_100000_M4 0.015

* ============================================================================
* Layer M5 - 12x12 grid
* ============================================================================

* M5 Horizontal resistors
r 8000_8000_M5 16000_8000_M5 0.010
r 16000_8000_M5 24000_8000_M5 0.010
r 24000_8000_M5 32000_8000_M5 0.010
r 32000_8000_M5 40000_8000_M5 0.010
r 40000_8000_M5 48000_8000_M5 0.010
r 48000_8000_M5 56000_8000_M5 0.010
r 56000_8000_M5 64000_8000_M5 0.010
r 64000_8000_M5 72000_8000_M5 0.010
r 72000_8000_M5 80000_8000_M5 0.010
r 80000_8000_M5 88000_8000_M5 0.010
r 88000_8000_M5 96000_8000_M5 0.010
r 8000_16000_M5 16000_16000_M5 0.010
r 16000_16000_M5 24000_16000_M5 0.010
r 24000_16000_M5 32000_16000_M5 0.010
r 32000_16000_M5 40000_16000_M5 0.010
r 40000_16000_M5 48000_16000_M5 0.010
r 48000_16000_M5 56000_16000_M5 0.010
r 56000_16000_M5 64000_16000_M5 0.010
r 64000_16000_M5 72000_16000_M5 0.010
r 72000_16000_M5 80000_16000_M5 0.010
r 80000_16000_M5 88000_16000_M5 0.010
r 88000_16000_M5 96000_16000_M5 0.010
r 8000_24000_M5 16000_24000_M5 0.010
r 16000_24000_M5 24000_24000_M5 0.010
r 24000_24000_M5 32000_24000_M5 0.010
r 32000_24000_M5 40000_24000_M5 0.010
r 40000_24000_M5 48000_24000_M5 0.010
r 48000_24000_M5 56000_24000_M5 0.010
r 56000_24000_M5 64000_24000_M5 0.010
r 64000_24000_M5 72000_24000_M5 0.010
r 72000_24000_M5 80000_24000_M5 0.010
r 80000_24000_M5 88000_24000_M5 0.010
r 88000_24000_M5 96000_24000_M5 0.010
r 8000_32000_M5 16000_32000_M5 0.010
r 16000_32000_M5 24000_32000_M5 0.010
r 24000_32000_M5 32000_32000_M5 0.010
r 32000_32000_M5 40000_32000_M5 0.010
r 40000_32000_M5 48000_32000_M5 0.010
r 48000_32000_M5 56000_32000_M5 0.010
r 56000_32000_M5 64000_32000_M5 0.010
r 64000_32000_M5 72000_32000_M5 0.010
r 72000_32000_M5 80000_32000_M5 0.010
r 80000_32000_M5 88000_32000_M5 0.010
r 88000_32000_M5 96000_32000_M5 0.010
r 8000_40000_M5 16000_40000_M5 0.010
r 16000_40000_M5 24000_40000_M5 0.010
r 24000_40000_M5 32000_40000_M5 0.010
r 32000_40000_M5 40000_40000_M5 0.010
r 40000_40000_M5 48000_40000_M5 0.010
r 48000_40000_M5 56000_40000_M5 0.010
r 56000_40000_M5 64000_40000_M5 0.010
r 64000_40000_M5 72000_40000_M5 0.010
r 72000_40000_M5 80000_40000_M5 0.010
r 80000_40000_M5 88000_40000_M5 0.010
r 88000_40000_M5 96000_40000_M5 0.010
r 8000_48000_M5 16000_48000_M5 0.010
r 16000_48000_M5 24000_48000_M5 0.010
r 24000_48000_M5 32000_48000_M5 0.010
r 32000_48000_M5 40000_48000_M5 0.010
r 40000_48000_M5 48000_48000_M5 0.010
r 48000_48000_M5 56000_48000_M5 0.010
r 56000_48000_M5 64000_48000_M5 0.010
r 64000_48000_M5 72000_48000_M5 0.010
r 72000_48000_M5 80000_48000_M5 0.010
r 80000_48000_M5 88000_48000_M5 0.010
r 88000_48000_M5 96000_48000_M5 0.010
r 8000_56000_M5 16000_56000_M5 0.010
r 16000_56000_M5 24000_56000_M5 0.010
r 24000_56000_M5 32000_56000_M5 0.010
r 32000_56000_M5 40000_56000_M5 0.010
r 40000_56000_M5 48000_56000_M5 0.010
r 48000_56000_M5 56000_56000_M5 0.010
r 56000_56000_M5 64000_56000_M5 0.010
r 64000_56000_M5 72000_56000_M5 0.010
r 72000_56000_M5 80000_56000_M5 0.010
r 80000_56000_M5 88000_56000_M5 0.010
r 88000_56000_M5 96000_56000_M5 0.010
r 8000_64000_M5 16000_64000_M5 0.010
r 16000_64000_M5 24000_64000_M5 0.010
r 24000_64000_M5 32000_64000_M5 0.010
r 32000_64000_M5 40000_64000_M5 0.010
r 40000_64000_M5 48000_64000_M5 0.010
r 48000_64000_M5 56000_64000_M5 0.010
r 56000_64000_M5 64000_64000_M5 0.010
r 64000_64000_M5 72000_64000_M5 0.010
r 72000_64000_M5 80000_64000_M5 0.010
r 80000_64000_M5 88000_64000_M5 0.010
r 88000_64000_M5 96000_64000_M5 0.010
r 8000_72000_M5 16000_72000_M5 0.010
r 16000_72000_M5 24000_72000_M5 0.010
r 24000_72000_M5 32000_72000_M5 0.010
r 32000_72000_M5 40000_72000_M5 0.010
r 40000_72000_M5 48000_72000_M5 0.010
r 48000_72000_M5 56000_72000_M5 0.010
r 56000_72000_M5 64000_72000_M5 0.010
r 64000_72000_M5 72000_72000_M5 0.010
r 72000_72000_M5 80000_72000_M5 0.010
r 80000_72000_M5 88000_72000_M5 0.010
r 88000_72000_M5 96000_72000_M5 0.010
r 8000_80000_M5 16000_80000_M5 0.010
r 16000_80000_M5 24000_80000_M5 0.010
r 24000_80000_M5 32000_80000_M5 0.010
r 32000_80000_M5 40000_80000_M5 0.010
r 40000_80000_M5 48000_80000_M5 0.010
r 48000_80000_M5 56000_80000_M5 0.010
r 56000_80000_M5 64000_80000_M5 0.010
r 64000_80000_M5 72000_80000_M5 0.010
r 72000_80000_M5 80000_80000_M5 0.010
r 80000_80000_M5 88000_80000_M5 0.010
r 88000_80000_M5 96000_80000_M5 0.010
r 8000_88000_M5 16000_88000_M5 0.010
r 16000_88000_M5 24000_88000_M5 0.010
r 24000_88000_M5 32000_88000_M5 0.010
r 32000_88000_M5 40000_88000_M5 0.010
r 40000_88000_M5 48000_88000_M5 0.010
r 48000_88000_M5 56000_88000_M5 0.010
r 56000_88000_M5 64000_88000_M5 0.010
r 64000_88000_M5 72000_88000_M5 0.010
r 72000_88000_M5 80000_88000_M5 0.010
r 80000_88000_M5 88000_88000_M5 0.010
r 88000_88000_M5 96000_88000_M5 0.010
r 8000_96000_M5 16000_96000_M5 0.010
r 16000_96000_M5 24000_96000_M5 0.010
r 24000_96000_M5 32000_96000_M5 0.010
r 32000_96000_M5 40000_96000_M5 0.010
r 40000_96000_M5 48000_96000_M5 0.010
r 48000_96000_M5 56000_96000_M5 0.010
r 56000_96000_M5 64000_96000_M5 0.010
r 64000_96000_M5 72000_96000_M5 0.010
r 72000_96000_M5 80000_96000_M5 0.010
r 80000_96000_M5 88000_96000_M5 0.010
r 88000_96000_M5 96000_96000_M5 0.010

* M5 Vertical resistors
r 8000_8000_M5 8000_16000_M5 0.012
r 8000_16000_M5 8000_24000_M5 0.012
r 8000_24000_M5 8000_32000_M5 0.012
r 8000_32000_M5 8000_40000_M5 0.012
r 8000_40000_M5 8000_48000_M5 0.012
r 8000_48000_M5 8000_56000_M5 0.012
r 8000_56000_M5 8000_64000_M5 0.012
r 8000_64000_M5 8000_72000_M5 0.012
r 8000_72000_M5 8000_80000_M5 0.012
r 8000_80000_M5 8000_88000_M5 0.012
r 8000_88000_M5 8000_96000_M5 0.012
r 16000_8000_M5 16000_16000_M5 0.012
r 16000_16000_M5 16000_24000_M5 0.012
r 16000_24000_M5 16000_32000_M5 0.012
r 16000_32000_M5 16000_40000_M5 0.012
r 16000_40000_M5 16000_48000_M5 0.012
r 16000_48000_M5 16000_56000_M5 0.012
r 16000_56000_M5 16000_64000_M5 0.012
r 16000_64000_M5 16000_72000_M5 0.012
r 16000_72000_M5 16000_80000_M5 0.012
r 16000_80000_M5 16000_88000_M5 0.012
r 16000_88000_M5 16000_96000_M5 0.012
r 24000_8000_M5 24000_16000_M5 0.012
r 24000_16000_M5 24000_24000_M5 0.012
r 24000_24000_M5 24000_32000_M5 0.012
r 24000_32000_M5 24000_40000_M5 0.012
r 24000_40000_M5 24000_48000_M5 0.012
r 24000_48000_M5 24000_56000_M5 0.012
r 24000_56000_M5 24000_64000_M5 0.012
r 24000_64000_M5 24000_72000_M5 0.012
r 24000_72000_M5 24000_80000_M5 0.012
r 24000_80000_M5 24000_88000_M5 0.012
r 24000_88000_M5 24000_96000_M5 0.012
r 32000_8000_M5 32000_16000_M5 0.012
r 32000_16000_M5 32000_24000_M5 0.012
r 32000_24000_M5 32000_32000_M5 0.012
r 32000_32000_M5 32000_40000_M5 0.012
r 32000_40000_M5 32000_48000_M5 0.012
r 32000_48000_M5 32000_56000_M5 0.012
r 32000_56000_M5 32000_64000_M5 0.012
r 32000_64000_M5 32000_72000_M5 0.012
r 32000_72000_M5 32000_80000_M5 0.012
r 32000_80000_M5 32000_88000_M5 0.012
r 32000_88000_M5 32000_96000_M5 0.012
r 40000_8000_M5 40000_16000_M5 0.012
r 40000_16000_M5 40000_24000_M5 0.012
r 40000_24000_M5 40000_32000_M5 0.012
r 40000_32000_M5 40000_40000_M5 0.012
r 40000_40000_M5 40000_48000_M5 0.012
r 40000_48000_M5 40000_56000_M5 0.012
r 40000_56000_M5 40000_64000_M5 0.012
r 40000_64000_M5 40000_72000_M5 0.012
r 40000_72000_M5 40000_80000_M5 0.012
r 40000_80000_M5 40000_88000_M5 0.012
r 40000_88000_M5 40000_96000_M5 0.012
r 48000_8000_M5 48000_16000_M5 0.012
r 48000_16000_M5 48000_24000_M5 0.012
r 48000_24000_M5 48000_32000_M5 0.012
r 48000_32000_M5 48000_40000_M5 0.012
r 48000_40000_M5 48000_48000_M5 0.012
r 48000_48000_M5 48000_56000_M5 0.012
r 48000_56000_M5 48000_64000_M5 0.012
r 48000_64000_M5 48000_72000_M5 0.012
r 48000_72000_M5 48000_80000_M5 0.012
r 48000_80000_M5 48000_88000_M5 0.012
r 48000_88000_M5 48000_96000_M5 0.012
r 56000_8000_M5 56000_16000_M5 0.012
r 56000_16000_M5 56000_24000_M5 0.012
r 56000_24000_M5 56000_32000_M5 0.012
r 56000_32000_M5 56000_40000_M5 0.012
r 56000_40000_M5 56000_48000_M5 0.012
r 56000_48000_M5 56000_56000_M5 0.012
r 56000_56000_M5 56000_64000_M5 0.012
r 56000_64000_M5 56000_72000_M5 0.012
r 56000_72000_M5 56000_80000_M5 0.012
r 56000_80000_M5 56000_88000_M5 0.012
r 56000_88000_M5 56000_96000_M5 0.012
r 64000_8000_M5 64000_16000_M5 0.012
r 64000_16000_M5 64000_24000_M5 0.012
r 64000_24000_M5 64000_32000_M5 0.012
r 64000_32000_M5 64000_40000_M5 0.012
r 64000_40000_M5 64000_48000_M5 0.012
r 64000_48000_M5 64000_56000_M5 0.012
r 64000_56000_M5 64000_64000_M5 0.012
r 64000_64000_M5 64000_72000_M5 0.012
r 64000_72000_M5 64000_80000_M5 0.012
r 64000_80000_M5 64000_88000_M5 0.012
r 64000_88000_M5 64000_96000_M5 0.012
r 72000_8000_M5 72000_16000_M5 0.012
r 72000_16000_M5 72000_24000_M5 0.012
r 72000_24000_M5 72000_32000_M5 0.012
r 72000_32000_M5 72000_40000_M5 0.012
r 72000_40000_M5 72000_48000_M5 0.012
r 72000_48000_M5 72000_56000_M5 0.012
r 72000_56000_M5 72000_64000_M5 0.012
r 72000_64000_M5 72000_72000_M5 0.012
r 72000_72000_M5 72000_80000_M5 0.012
r 72000_80000_M5 72000_88000_M5 0.012
r 72000_88000_M5 72000_96000_M5 0.012
r 80000_8000_M5 80000_16000_M5 0.012
r 80000_16000_M5 80000_24000_M5 0.012
r 80000_24000_M5 80000_32000_M5 0.012
r 80000_32000_M5 80000_40000_M5 0.012
r 80000_40000_M5 80000_48000_M5 0.012
r 80000_48000_M5 80000_56000_M5 0.012
r 80000_56000_M5 80000_64000_M5 0.012
r 80000_64000_M5 80000_72000_M5 0.012
r 80000_72000_M5 80000_80000_M5 0.012
r 80000_80000_M5 80000_88000_M5 0.012
r 80000_88000_M5 80000_96000_M5 0.012
r 88000_8000_M5 88000_16000_M5 0.012
r 88000_16000_M5 88000_24000_M5 0.012
r 88000_24000_M5 88000_32000_M5 0.012
r 88000_32000_M5 88000_40000_M5 0.012
r 88000_40000_M5 88000_48000_M5 0.012
r 88000_48000_M5 88000_56000_M5 0.012
r 88000_56000_M5 88000_64000_M5 0.012
r 88000_64000_M5 88000_72000_M5 0.012
r 88000_72000_M5 88000_80000_M5 0.012
r 88000_80000_M5 88000_88000_M5 0.012
r 88000_88000_M5 88000_96000_M5 0.012
r 96000_8000_M5 96000_16000_M5 0.012
r 96000_16000_M5 96000_24000_M5 0.012
r 96000_24000_M5 96000_32000_M5 0.012
r 96000_32000_M5 96000_40000_M5 0.012
r 96000_40000_M5 96000_48000_M5 0.012
r 96000_48000_M5 96000_56000_M5 0.012
r 96000_56000_M5 96000_64000_M5 0.012
r 96000_64000_M5 96000_72000_M5 0.012
r 96000_72000_M5 96000_80000_M5 0.012
r 96000_80000_M5 96000_88000_M5 0.012
r 96000_88000_M5 96000_96000_M5 0.012

* ============================================================================
* Via connections M1 to M2
* ============================================================================

r 2000_2000_M1 2000_2000_M2 0.050
r 2000_4000_M1 2000_4000_M2 0.050
r 2000_6000_M1 2000_6000_M2 0.050
r 2000_8000_M1 2000_8000_M2 0.050
r 2000_10000_M1 2000_10000_M2 0.050
r 2000_12000_M1 2000_12000_M2 0.050
r 2000_14000_M1 2000_14000_M2 0.050
r 2000_16000_M1 2000_16000_M2 0.050
r 2000_18000_M1 2000_18000_M2 0.050
r 2000_20000_M1 2000_20000_M2 0.050
r 2000_22000_M1 2000_22000_M2 0.050
r 2000_24000_M1 2000_24000_M2 0.050
r 2000_26000_M1 2000_26000_M2 0.050
r 2000_28000_M1 2000_28000_M2 0.050
r 2000_30000_M1 2000_30000_M2 0.050
r 2000_32000_M1 2000_32000_M2 0.050
r 2000_34000_M1 2000_34000_M2 0.050
r 2000_36000_M1 2000_36000_M2 0.050
r 2000_38000_M1 2000_38000_M2 0.050
r 2000_40000_M1 2000_40000_M2 0.050
r 2000_42000_M1 2000_42000_M2 0.050
r 2000_44000_M1 2000_44000_M2 0.050
r 2000_46000_M1 2000_46000_M2 0.050
r 2000_48000_M1 2000_48000_M2 0.050
r 2000_50000_M1 2000_50000_M2 0.050
r 2000_52000_M1 2000_52000_M2 0.050
r 2000_54000_M1 2000_54000_M2 0.050
r 2000_56000_M1 2000_56000_M2 0.050
r 2000_58000_M1 2000_58000_M2 0.050
r 2000_60000_M1 2000_60000_M2 0.050
r 2000_62000_M1 2000_62000_M2 0.050
r 2000_64000_M1 2000_64000_M2 0.050
r 2000_66000_M1 2000_66000_M2 0.050
r 2000_68000_M1 2000_68000_M2 0.050
r 2000_70000_M1 2000_70000_M2 0.050
r 2000_72000_M1 2000_72000_M2 0.050
r 2000_74000_M1 2000_74000_M2 0.050
r 2000_76000_M1 2000_76000_M2 0.050
r 2000_78000_M1 2000_78000_M2 0.050
r 2000_80000_M1 2000_80000_M2 0.050
r 2000_82000_M1 2000_82000_M2 0.050
r 2000_84000_M1 2000_84000_M2 0.050
r 2000_86000_M1 2000_86000_M2 0.050
r 2000_88000_M1 2000_88000_M2 0.050
r 2000_90000_M1 2000_90000_M2 0.050
r 2000_92000_M1 2000_92000_M2 0.050
r 2000_94000_M1 2000_94000_M2 0.050
r 2000_96000_M1 2000_96000_M2 0.050
r 2000_98000_M1 2000_98000_M2 0.050
r 2000_100000_M1 2000_100000_M2 0.050
r 4000_2000_M1 4000_2000_M2 0.050
r 4000_4000_M1 4000_4000_M2 0.050
r 4000_6000_M1 4000_6000_M2 0.050
r 4000_8000_M1 4000_8000_M2 0.050
r 4000_10000_M1 4000_10000_M2 0.050
r 4000_12000_M1 4000_12000_M2 0.050
r 4000_14000_M1 4000_14000_M2 0.050
r 4000_16000_M1 4000_16000_M2 0.050
r 4000_18000_M1 4000_18000_M2 0.050
r 4000_20000_M1 4000_20000_M2 0.050
r 4000_22000_M1 4000_22000_M2 0.050
r 4000_24000_M1 4000_24000_M2 0.050
r 4000_26000_M1 4000_26000_M2 0.050
r 4000_28000_M1 4000_28000_M2 0.050
r 4000_30000_M1 4000_30000_M2 0.050
r 4000_32000_M1 4000_32000_M2 0.050
r 4000_34000_M1 4000_34000_M2 0.050
r 4000_36000_M1 4000_36000_M2 0.050
r 4000_38000_M1 4000_38000_M2 0.050
r 4000_40000_M1 4000_40000_M2 0.050
r 4000_42000_M1 4000_42000_M2 0.050
r 4000_44000_M1 4000_44000_M2 0.050
r 4000_46000_M1 4000_46000_M2 0.050
r 4000_48000_M1 4000_48000_M2 0.050
r 4000_50000_M1 4000_50000_M2 0.050
r 4000_52000_M1 4000_52000_M2 0.050
r 4000_54000_M1 4000_54000_M2 0.050
r 4000_56000_M1 4000_56000_M2 0.050
r 4000_58000_M1 4000_58000_M2 0.050
r 4000_60000_M1 4000_60000_M2 0.050
r 4000_62000_M1 4000_62000_M2 0.050
r 4000_64000_M1 4000_64000_M2 0.050
r 4000_66000_M1 4000_66000_M2 0.050
r 4000_68000_M1 4000_68000_M2 0.050
r 4000_70000_M1 4000_70000_M2 0.050
r 4000_72000_M1 4000_72000_M2 0.050
r 4000_74000_M1 4000_74000_M2 0.050
r 4000_76000_M1 4000_76000_M2 0.050
r 4000_78000_M1 4000_78000_M2 0.050
r 4000_80000_M1 4000_80000_M2 0.050
r 4000_82000_M1 4000_82000_M2 0.050
r 4000_84000_M1 4000_84000_M2 0.050
r 4000_86000_M1 4000_86000_M2 0.050
r 4000_88000_M1 4000_88000_M2 0.050
r 4000_90000_M1 4000_90000_M2 0.050
r 4000_92000_M1 4000_92000_M2 0.050
r 4000_94000_M1 4000_94000_M2 0.050
r 4000_96000_M1 4000_96000_M2 0.050
r 4000_98000_M1 4000_98000_M2 0.050
r 4000_100000_M1 4000_100000_M2 0.050
r 6000_2000_M1 6000_2000_M2 0.050
r 6000_4000_M1 6000_4000_M2 0.050
r 6000_6000_M1 6000_6000_M2 0.050
r 6000_8000_M1 6000_8000_M2 0.050
r 6000_10000_M1 6000_10000_M2 0.050
r 6000_12000_M1 6000_12000_M2 0.050
r 6000_14000_M1 6000_14000_M2 0.050
r 6000_16000_M1 6000_16000_M2 0.050
r 6000_18000_M1 6000_18000_M2 0.050
r 6000_20000_M1 6000_20000_M2 0.050
r 6000_22000_M1 6000_22000_M2 0.050
r 6000_24000_M1 6000_24000_M2 0.050
r 6000_26000_M1 6000_26000_M2 0.050
r 6000_28000_M1 6000_28000_M2 0.050
r 6000_30000_M1 6000_30000_M2 0.050
r 6000_32000_M1 6000_32000_M2 0.050
r 6000_34000_M1 6000_34000_M2 0.050
r 6000_36000_M1 6000_36000_M2 0.050
r 6000_38000_M1 6000_38000_M2 0.050
r 6000_40000_M1 6000_40000_M2 0.050
r 6000_42000_M1 6000_42000_M2 0.050
r 6000_44000_M1 6000_44000_M2 0.050
r 6000_46000_M1 6000_46000_M2 0.050
r 6000_48000_M1 6000_48000_M2 0.050
r 6000_50000_M1 6000_50000_M2 0.050
r 6000_52000_M1 6000_52000_M2 0.050
r 6000_54000_M1 6000_54000_M2 0.050
r 6000_56000_M1 6000_56000_M2 0.050
r 6000_58000_M1 6000_58000_M2 0.050
r 6000_60000_M1 6000_60000_M2 0.050
r 6000_62000_M1 6000_62000_M2 0.050
r 6000_64000_M1 6000_64000_M2 0.050
r 6000_66000_M1 6000_66000_M2 0.050
r 6000_68000_M1 6000_68000_M2 0.050
r 6000_70000_M1 6000_70000_M2 0.050
r 6000_72000_M1 6000_72000_M2 0.050
r 6000_74000_M1 6000_74000_M2 0.050
r 6000_76000_M1 6000_76000_M2 0.050
r 6000_78000_M1 6000_78000_M2 0.050
r 6000_80000_M1 6000_80000_M2 0.050
r 6000_82000_M1 6000_82000_M2 0.050
r 6000_84000_M1 6000_84000_M2 0.050
r 6000_86000_M1 6000_86000_M2 0.050
r 6000_88000_M1 6000_88000_M2 0.050
r 6000_90000_M1 6000_90000_M2 0.050
r 6000_92000_M1 6000_92000_M2 0.050
r 6000_94000_M1 6000_94000_M2 0.050
r 6000_96000_M1 6000_96000_M2 0.050
r 6000_98000_M1 6000_98000_M2 0.050
r 6000_100000_M1 6000_100000_M2 0.050
r 8000_2000_M1 8000_2000_M2 0.050
r 8000_4000_M1 8000_4000_M2 0.050
r 8000_6000_M1 8000_6000_M2 0.050
r 8000_8000_M1 8000_8000_M2 0.050
r 8000_10000_M1 8000_10000_M2 0.050
r 8000_12000_M1 8000_12000_M2 0.050
r 8000_14000_M1 8000_14000_M2 0.050
r 8000_16000_M1 8000_16000_M2 0.050
r 8000_18000_M1 8000_18000_M2 0.050
r 8000_20000_M1 8000_20000_M2 0.050
r 8000_22000_M1 8000_22000_M2 0.050
r 8000_24000_M1 8000_24000_M2 0.050
r 8000_26000_M1 8000_26000_M2 0.050
r 8000_28000_M1 8000_28000_M2 0.050
r 8000_30000_M1 8000_30000_M2 0.050
r 8000_32000_M1 8000_32000_M2 0.050
r 8000_34000_M1 8000_34000_M2 0.050
r 8000_36000_M1 8000_36000_M2 0.050
r 8000_38000_M1 8000_38000_M2 0.050
r 8000_40000_M1 8000_40000_M2 0.050
r 8000_42000_M1 8000_42000_M2 0.050
r 8000_44000_M1 8000_44000_M2 0.050
r 8000_46000_M1 8000_46000_M2 0.050
r 8000_48000_M1 8000_48000_M2 0.050
r 8000_50000_M1 8000_50000_M2 0.050
r 8000_52000_M1 8000_52000_M2 0.050
r 8000_54000_M1 8000_54000_M2 0.050
r 8000_56000_M1 8000_56000_M2 0.050
r 8000_58000_M1 8000_58000_M2 0.050
r 8000_60000_M1 8000_60000_M2 0.050
r 8000_62000_M1 8000_62000_M2 0.050
r 8000_64000_M1 8000_64000_M2 0.050
r 8000_66000_M1 8000_66000_M2 0.050
r 8000_68000_M1 8000_68000_M2 0.050
r 8000_70000_M1 8000_70000_M2 0.050
r 8000_72000_M1 8000_72000_M2 0.050
r 8000_74000_M1 8000_74000_M2 0.050
r 8000_76000_M1 8000_76000_M2 0.050
r 8000_78000_M1 8000_78000_M2 0.050
r 8000_80000_M1 8000_80000_M2 0.050
r 8000_82000_M1 8000_82000_M2 0.050
r 8000_84000_M1 8000_84000_M2 0.050
r 8000_86000_M1 8000_86000_M2 0.050
r 8000_88000_M1 8000_88000_M2 0.050
r 8000_90000_M1 8000_90000_M2 0.050
r 8000_92000_M1 8000_92000_M2 0.050
r 8000_94000_M1 8000_94000_M2 0.050
r 8000_96000_M1 8000_96000_M2 0.050
r 8000_98000_M1 8000_98000_M2 0.050
r 8000_100000_M1 8000_100000_M2 0.050
r 10000_2000_M1 10000_2000_M2 0.050
r 10000_4000_M1 10000_4000_M2 0.050
r 10000_6000_M1 10000_6000_M2 0.050
r 10000_8000_M1 10000_8000_M2 0.050
r 10000_10000_M1 10000_10000_M2 0.050
r 10000_12000_M1 10000_12000_M2 0.050
r 10000_14000_M1 10000_14000_M2 0.050
r 10000_16000_M1 10000_16000_M2 0.050
r 10000_18000_M1 10000_18000_M2 0.050
r 10000_20000_M1 10000_20000_M2 0.050
r 10000_22000_M1 10000_22000_M2 0.050
r 10000_24000_M1 10000_24000_M2 0.050
r 10000_26000_M1 10000_26000_M2 0.050
r 10000_28000_M1 10000_28000_M2 0.050
r 10000_30000_M1 10000_30000_M2 0.050
r 10000_32000_M1 10000_32000_M2 0.050
r 10000_34000_M1 10000_34000_M2 0.050
r 10000_36000_M1 10000_36000_M2 0.050
r 10000_38000_M1 10000_38000_M2 0.050
r 10000_40000_M1 10000_40000_M2 0.050
r 10000_42000_M1 10000_42000_M2 0.050
r 10000_44000_M1 10000_44000_M2 0.050
r 10000_46000_M1 10000_46000_M2 0.050
r 10000_48000_M1 10000_48000_M2 0.050
r 10000_50000_M1 10000_50000_M2 0.050
r 10000_52000_M1 10000_52000_M2 0.050
r 10000_54000_M1 10000_54000_M2 0.050
r 10000_56000_M1 10000_56000_M2 0.050
r 10000_58000_M1 10000_58000_M2 0.050
r 10000_60000_M1 10000_60000_M2 0.050
r 10000_62000_M1 10000_62000_M2 0.050
r 10000_64000_M1 10000_64000_M2 0.050
r 10000_66000_M1 10000_66000_M2 0.050
r 10000_68000_M1 10000_68000_M2 0.050
r 10000_70000_M1 10000_70000_M2 0.050
r 10000_72000_M1 10000_72000_M2 0.050
r 10000_74000_M1 10000_74000_M2 0.050
r 10000_76000_M1 10000_76000_M2 0.050
r 10000_78000_M1 10000_78000_M2 0.050
r 10000_80000_M1 10000_80000_M2 0.050
r 10000_82000_M1 10000_82000_M2 0.050
r 10000_84000_M1 10000_84000_M2 0.050
r 10000_86000_M1 10000_86000_M2 0.050
r 10000_88000_M1 10000_88000_M2 0.050
r 10000_90000_M1 10000_90000_M2 0.050
r 10000_92000_M1 10000_92000_M2 0.050
r 10000_94000_M1 10000_94000_M2 0.050
r 10000_96000_M1 10000_96000_M2 0.050
r 10000_98000_M1 10000_98000_M2 0.050
r 10000_100000_M1 10000_100000_M2 0.050
r 12000_2000_M1 12000_2000_M2 0.050
r 12000_4000_M1 12000_4000_M2 0.050
r 12000_6000_M1 12000_6000_M2 0.050
r 12000_8000_M1 12000_8000_M2 0.050
r 12000_10000_M1 12000_10000_M2 0.050
r 12000_12000_M1 12000_12000_M2 0.050
r 12000_14000_M1 12000_14000_M2 0.050
r 12000_16000_M1 12000_16000_M2 0.050
r 12000_18000_M1 12000_18000_M2 0.050
r 12000_20000_M1 12000_20000_M2 0.050
r 12000_22000_M1 12000_22000_M2 0.050
r 12000_24000_M1 12000_24000_M2 0.050
r 12000_26000_M1 12000_26000_M2 0.050
r 12000_28000_M1 12000_28000_M2 0.050
r 12000_30000_M1 12000_30000_M2 0.050
r 12000_32000_M1 12000_32000_M2 0.050
r 12000_34000_M1 12000_34000_M2 0.050
r 12000_36000_M1 12000_36000_M2 0.050
r 12000_38000_M1 12000_38000_M2 0.050
r 12000_40000_M1 12000_40000_M2 0.050
r 12000_42000_M1 12000_42000_M2 0.050
r 12000_44000_M1 12000_44000_M2 0.050
r 12000_46000_M1 12000_46000_M2 0.050
r 12000_48000_M1 12000_48000_M2 0.050
r 12000_50000_M1 12000_50000_M2 0.050
r 12000_52000_M1 12000_52000_M2 0.050
r 12000_54000_M1 12000_54000_M2 0.050
r 12000_56000_M1 12000_56000_M2 0.050
r 12000_58000_M1 12000_58000_M2 0.050
r 12000_60000_M1 12000_60000_M2 0.050
r 12000_62000_M1 12000_62000_M2 0.050
r 12000_64000_M1 12000_64000_M2 0.050
r 12000_66000_M1 12000_66000_M2 0.050
r 12000_68000_M1 12000_68000_M2 0.050
r 12000_70000_M1 12000_70000_M2 0.050
r 12000_72000_M1 12000_72000_M2 0.050
r 12000_74000_M1 12000_74000_M2 0.050
r 12000_76000_M1 12000_76000_M2 0.050
r 12000_78000_M1 12000_78000_M2 0.050
r 12000_80000_M1 12000_80000_M2 0.050
r 12000_82000_M1 12000_82000_M2 0.050
r 12000_84000_M1 12000_84000_M2 0.050
r 12000_86000_M1 12000_86000_M2 0.050
r 12000_88000_M1 12000_88000_M2 0.050
r 12000_90000_M1 12000_90000_M2 0.050
r 12000_92000_M1 12000_92000_M2 0.050
r 12000_94000_M1 12000_94000_M2 0.050
r 12000_96000_M1 12000_96000_M2 0.050
r 12000_98000_M1 12000_98000_M2 0.050
r 12000_100000_M1 12000_100000_M2 0.050
r 14000_2000_M1 14000_2000_M2 0.050
r 14000_4000_M1 14000_4000_M2 0.050
r 14000_6000_M1 14000_6000_M2 0.050
r 14000_8000_M1 14000_8000_M2 0.050
r 14000_10000_M1 14000_10000_M2 0.050
r 14000_12000_M1 14000_12000_M2 0.050
r 14000_14000_M1 14000_14000_M2 0.050
r 14000_16000_M1 14000_16000_M2 0.050
r 14000_18000_M1 14000_18000_M2 0.050
r 14000_20000_M1 14000_20000_M2 0.050
r 14000_22000_M1 14000_22000_M2 0.050
r 14000_24000_M1 14000_24000_M2 0.050
r 14000_26000_M1 14000_26000_M2 0.050
r 14000_28000_M1 14000_28000_M2 0.050
r 14000_30000_M1 14000_30000_M2 0.050
r 14000_32000_M1 14000_32000_M2 0.050
r 14000_34000_M1 14000_34000_M2 0.050
r 14000_36000_M1 14000_36000_M2 0.050
r 14000_38000_M1 14000_38000_M2 0.050
r 14000_40000_M1 14000_40000_M2 0.050
r 14000_42000_M1 14000_42000_M2 0.050
r 14000_44000_M1 14000_44000_M2 0.050
r 14000_46000_M1 14000_46000_M2 0.050
r 14000_48000_M1 14000_48000_M2 0.050
r 14000_50000_M1 14000_50000_M2 0.050
r 14000_52000_M1 14000_52000_M2 0.050
r 14000_54000_M1 14000_54000_M2 0.050
r 14000_56000_M1 14000_56000_M2 0.050
r 14000_58000_M1 14000_58000_M2 0.050
r 14000_60000_M1 14000_60000_M2 0.050
r 14000_62000_M1 14000_62000_M2 0.050
r 14000_64000_M1 14000_64000_M2 0.050
r 14000_66000_M1 14000_66000_M2 0.050
r 14000_68000_M1 14000_68000_M2 0.050
r 14000_70000_M1 14000_70000_M2 0.050
r 14000_72000_M1 14000_72000_M2 0.050
r 14000_74000_M1 14000_74000_M2 0.050
r 14000_76000_M1 14000_76000_M2 0.050
r 14000_78000_M1 14000_78000_M2 0.050
r 14000_80000_M1 14000_80000_M2 0.050
r 14000_82000_M1 14000_82000_M2 0.050
r 14000_84000_M1 14000_84000_M2 0.050
r 14000_86000_M1 14000_86000_M2 0.050
r 14000_88000_M1 14000_88000_M2 0.050
r 14000_90000_M1 14000_90000_M2 0.050
r 14000_92000_M1 14000_92000_M2 0.050
r 14000_94000_M1 14000_94000_M2 0.050
r 14000_96000_M1 14000_96000_M2 0.050
r 14000_98000_M1 14000_98000_M2 0.050
r 14000_100000_M1 14000_100000_M2 0.050
r 16000_2000_M1 16000_2000_M2 0.050
r 16000_4000_M1 16000_4000_M2 0.050
r 16000_6000_M1 16000_6000_M2 0.050
r 16000_8000_M1 16000_8000_M2 0.050
r 16000_10000_M1 16000_10000_M2 0.050
r 16000_12000_M1 16000_12000_M2 0.050
r 16000_14000_M1 16000_14000_M2 0.050
r 16000_16000_M1 16000_16000_M2 0.050
r 16000_18000_M1 16000_18000_M2 0.050
r 16000_20000_M1 16000_20000_M2 0.050
r 16000_22000_M1 16000_22000_M2 0.050
r 16000_24000_M1 16000_24000_M2 0.050
r 16000_26000_M1 16000_26000_M2 0.050
r 16000_28000_M1 16000_28000_M2 0.050
r 16000_30000_M1 16000_30000_M2 0.050
r 16000_32000_M1 16000_32000_M2 0.050
r 16000_34000_M1 16000_34000_M2 0.050
r 16000_36000_M1 16000_36000_M2 0.050
r 16000_38000_M1 16000_38000_M2 0.050
r 16000_40000_M1 16000_40000_M2 0.050
r 16000_42000_M1 16000_42000_M2 0.050
r 16000_44000_M1 16000_44000_M2 0.050
r 16000_46000_M1 16000_46000_M2 0.050
r 16000_48000_M1 16000_48000_M2 0.050
r 16000_50000_M1 16000_50000_M2 0.050
r 16000_52000_M1 16000_52000_M2 0.050
r 16000_54000_M1 16000_54000_M2 0.050
r 16000_56000_M1 16000_56000_M2 0.050
r 16000_58000_M1 16000_58000_M2 0.050
r 16000_60000_M1 16000_60000_M2 0.050
r 16000_62000_M1 16000_62000_M2 0.050
r 16000_64000_M1 16000_64000_M2 0.050
r 16000_66000_M1 16000_66000_M2 0.050
r 16000_68000_M1 16000_68000_M2 0.050
r 16000_70000_M1 16000_70000_M2 0.050
r 16000_72000_M1 16000_72000_M2 0.050
r 16000_74000_M1 16000_74000_M2 0.050
r 16000_76000_M1 16000_76000_M2 0.050
r 16000_78000_M1 16000_78000_M2 0.050
r 16000_80000_M1 16000_80000_M2 0.050
r 16000_82000_M1 16000_82000_M2 0.050
r 16000_84000_M1 16000_84000_M2 0.050
r 16000_86000_M1 16000_86000_M2 0.050
r 16000_88000_M1 16000_88000_M2 0.050
r 16000_90000_M1 16000_90000_M2 0.050
r 16000_92000_M1 16000_92000_M2 0.050
r 16000_94000_M1 16000_94000_M2 0.050
r 16000_96000_M1 16000_96000_M2 0.050
r 16000_98000_M1 16000_98000_M2 0.050
r 16000_100000_M1 16000_100000_M2 0.050
r 18000_2000_M1 18000_2000_M2 0.050
r 18000_4000_M1 18000_4000_M2 0.050
r 18000_6000_M1 18000_6000_M2 0.050
r 18000_8000_M1 18000_8000_M2 0.050
r 18000_10000_M1 18000_10000_M2 0.050
r 18000_12000_M1 18000_12000_M2 0.050
r 18000_14000_M1 18000_14000_M2 0.050
r 18000_16000_M1 18000_16000_M2 0.050
r 18000_18000_M1 18000_18000_M2 0.050
r 18000_20000_M1 18000_20000_M2 0.050
r 18000_22000_M1 18000_22000_M2 0.050
r 18000_24000_M1 18000_24000_M2 0.050
r 18000_26000_M1 18000_26000_M2 0.050
r 18000_28000_M1 18000_28000_M2 0.050
r 18000_30000_M1 18000_30000_M2 0.050
r 18000_32000_M1 18000_32000_M2 0.050
r 18000_34000_M1 18000_34000_M2 0.050
r 18000_36000_M1 18000_36000_M2 0.050
r 18000_38000_M1 18000_38000_M2 0.050
r 18000_40000_M1 18000_40000_M2 0.050
r 18000_42000_M1 18000_42000_M2 0.050
r 18000_44000_M1 18000_44000_M2 0.050
r 18000_46000_M1 18000_46000_M2 0.050
r 18000_48000_M1 18000_48000_M2 0.050
r 18000_50000_M1 18000_50000_M2 0.050
r 18000_52000_M1 18000_52000_M2 0.050
r 18000_54000_M1 18000_54000_M2 0.050
r 18000_56000_M1 18000_56000_M2 0.050
r 18000_58000_M1 18000_58000_M2 0.050
r 18000_60000_M1 18000_60000_M2 0.050
r 18000_62000_M1 18000_62000_M2 0.050
r 18000_64000_M1 18000_64000_M2 0.050
r 18000_66000_M1 18000_66000_M2 0.050
r 18000_68000_M1 18000_68000_M2 0.050
r 18000_70000_M1 18000_70000_M2 0.050
r 18000_72000_M1 18000_72000_M2 0.050
r 18000_74000_M1 18000_74000_M2 0.050
r 18000_76000_M1 18000_76000_M2 0.050
r 18000_78000_M1 18000_78000_M2 0.050
r 18000_80000_M1 18000_80000_M2 0.050
r 18000_82000_M1 18000_82000_M2 0.050
r 18000_84000_M1 18000_84000_M2 0.050
r 18000_86000_M1 18000_86000_M2 0.050
r 18000_88000_M1 18000_88000_M2 0.050
r 18000_90000_M1 18000_90000_M2 0.050
r 18000_92000_M1 18000_92000_M2 0.050
r 18000_94000_M1 18000_94000_M2 0.050
r 18000_96000_M1 18000_96000_M2 0.050
r 18000_98000_M1 18000_98000_M2 0.050
r 18000_100000_M1 18000_100000_M2 0.050
r 20000_2000_M1 20000_2000_M2 0.050
r 20000_4000_M1 20000_4000_M2 0.050
r 20000_6000_M1 20000_6000_M2 0.050
r 20000_8000_M1 20000_8000_M2 0.050
r 20000_10000_M1 20000_10000_M2 0.050
r 20000_12000_M1 20000_12000_M2 0.050
r 20000_14000_M1 20000_14000_M2 0.050
r 20000_16000_M1 20000_16000_M2 0.050
r 20000_18000_M1 20000_18000_M2 0.050
r 20000_20000_M1 20000_20000_M2 0.050
r 20000_22000_M1 20000_22000_M2 0.050
r 20000_24000_M1 20000_24000_M2 0.050
r 20000_26000_M1 20000_26000_M2 0.050
r 20000_28000_M1 20000_28000_M2 0.050
r 20000_30000_M1 20000_30000_M2 0.050
r 20000_32000_M1 20000_32000_M2 0.050
r 20000_34000_M1 20000_34000_M2 0.050
r 20000_36000_M1 20000_36000_M2 0.050
r 20000_38000_M1 20000_38000_M2 0.050
r 20000_40000_M1 20000_40000_M2 0.050
r 20000_42000_M1 20000_42000_M2 0.050
r 20000_44000_M1 20000_44000_M2 0.050
r 20000_46000_M1 20000_46000_M2 0.050
r 20000_48000_M1 20000_48000_M2 0.050
r 20000_50000_M1 20000_50000_M2 0.050
r 20000_52000_M1 20000_52000_M2 0.050
r 20000_54000_M1 20000_54000_M2 0.050
r 20000_56000_M1 20000_56000_M2 0.050
r 20000_58000_M1 20000_58000_M2 0.050
r 20000_60000_M1 20000_60000_M2 0.050
r 20000_62000_M1 20000_62000_M2 0.050
r 20000_64000_M1 20000_64000_M2 0.050
r 20000_66000_M1 20000_66000_M2 0.050
r 20000_68000_M1 20000_68000_M2 0.050
r 20000_70000_M1 20000_70000_M2 0.050
r 20000_72000_M1 20000_72000_M2 0.050
r 20000_74000_M1 20000_74000_M2 0.050
r 20000_76000_M1 20000_76000_M2 0.050
r 20000_78000_M1 20000_78000_M2 0.050
r 20000_80000_M1 20000_80000_M2 0.050
r 20000_82000_M1 20000_82000_M2 0.050
r 20000_84000_M1 20000_84000_M2 0.050
r 20000_86000_M1 20000_86000_M2 0.050
r 20000_88000_M1 20000_88000_M2 0.050
r 20000_90000_M1 20000_90000_M2 0.050
r 20000_92000_M1 20000_92000_M2 0.050
r 20000_94000_M1 20000_94000_M2 0.050
r 20000_96000_M1 20000_96000_M2 0.050
r 20000_98000_M1 20000_98000_M2 0.050
r 20000_100000_M1 20000_100000_M2 0.050
r 22000_2000_M1 22000_2000_M2 0.050
r 22000_4000_M1 22000_4000_M2 0.050
r 22000_6000_M1 22000_6000_M2 0.050
r 22000_8000_M1 22000_8000_M2 0.050
r 22000_10000_M1 22000_10000_M2 0.050
r 22000_12000_M1 22000_12000_M2 0.050
r 22000_14000_M1 22000_14000_M2 0.050
r 22000_16000_M1 22000_16000_M2 0.050
r 22000_18000_M1 22000_18000_M2 0.050
r 22000_20000_M1 22000_20000_M2 0.050
r 22000_22000_M1 22000_22000_M2 0.050
r 22000_24000_M1 22000_24000_M2 0.050
r 22000_26000_M1 22000_26000_M2 0.050
r 22000_28000_M1 22000_28000_M2 0.050
r 22000_30000_M1 22000_30000_M2 0.050
r 22000_32000_M1 22000_32000_M2 0.050
r 22000_34000_M1 22000_34000_M2 0.050
r 22000_36000_M1 22000_36000_M2 0.050
r 22000_38000_M1 22000_38000_M2 0.050
r 22000_40000_M1 22000_40000_M2 0.050
r 22000_42000_M1 22000_42000_M2 0.050
r 22000_44000_M1 22000_44000_M2 0.050
r 22000_46000_M1 22000_46000_M2 0.050
r 22000_48000_M1 22000_48000_M2 0.050
r 22000_50000_M1 22000_50000_M2 0.050
r 22000_52000_M1 22000_52000_M2 0.050
r 22000_54000_M1 22000_54000_M2 0.050
r 22000_56000_M1 22000_56000_M2 0.050
r 22000_58000_M1 22000_58000_M2 0.050
r 22000_60000_M1 22000_60000_M2 0.050
r 22000_62000_M1 22000_62000_M2 0.050
r 22000_64000_M1 22000_64000_M2 0.050
r 22000_66000_M1 22000_66000_M2 0.050
r 22000_68000_M1 22000_68000_M2 0.050
r 22000_70000_M1 22000_70000_M2 0.050
r 22000_72000_M1 22000_72000_M2 0.050
r 22000_74000_M1 22000_74000_M2 0.050
r 22000_76000_M1 22000_76000_M2 0.050
r 22000_78000_M1 22000_78000_M2 0.050
r 22000_80000_M1 22000_80000_M2 0.050
r 22000_82000_M1 22000_82000_M2 0.050
r 22000_84000_M1 22000_84000_M2 0.050
r 22000_86000_M1 22000_86000_M2 0.050
r 22000_88000_M1 22000_88000_M2 0.050
r 22000_90000_M1 22000_90000_M2 0.050
r 22000_92000_M1 22000_92000_M2 0.050
r 22000_94000_M1 22000_94000_M2 0.050
r 22000_96000_M1 22000_96000_M2 0.050
r 22000_98000_M1 22000_98000_M2 0.050
r 22000_100000_M1 22000_100000_M2 0.050
r 24000_2000_M1 24000_2000_M2 0.050
r 24000_4000_M1 24000_4000_M2 0.050
r 24000_6000_M1 24000_6000_M2 0.050
r 24000_8000_M1 24000_8000_M2 0.050
r 24000_10000_M1 24000_10000_M2 0.050
r 24000_12000_M1 24000_12000_M2 0.050
r 24000_14000_M1 24000_14000_M2 0.050
r 24000_16000_M1 24000_16000_M2 0.050
r 24000_18000_M1 24000_18000_M2 0.050
r 24000_20000_M1 24000_20000_M2 0.050
r 24000_22000_M1 24000_22000_M2 0.050
r 24000_24000_M1 24000_24000_M2 0.050
r 24000_26000_M1 24000_26000_M2 0.050
r 24000_28000_M1 24000_28000_M2 0.050
r 24000_30000_M1 24000_30000_M2 0.050
r 24000_32000_M1 24000_32000_M2 0.050
r 24000_34000_M1 24000_34000_M2 0.050
r 24000_36000_M1 24000_36000_M2 0.050
r 24000_38000_M1 24000_38000_M2 0.050
r 24000_40000_M1 24000_40000_M2 0.050
r 24000_42000_M1 24000_42000_M2 0.050
r 24000_44000_M1 24000_44000_M2 0.050
r 24000_46000_M1 24000_46000_M2 0.050
r 24000_48000_M1 24000_48000_M2 0.050
r 24000_50000_M1 24000_50000_M2 0.050
r 24000_52000_M1 24000_52000_M2 0.050
r 24000_54000_M1 24000_54000_M2 0.050
r 24000_56000_M1 24000_56000_M2 0.050
r 24000_58000_M1 24000_58000_M2 0.050
r 24000_60000_M1 24000_60000_M2 0.050
r 24000_62000_M1 24000_62000_M2 0.050
r 24000_64000_M1 24000_64000_M2 0.050
r 24000_66000_M1 24000_66000_M2 0.050
r 24000_68000_M1 24000_68000_M2 0.050
r 24000_70000_M1 24000_70000_M2 0.050
r 24000_72000_M1 24000_72000_M2 0.050
r 24000_74000_M1 24000_74000_M2 0.050
r 24000_76000_M1 24000_76000_M2 0.050
r 24000_78000_M1 24000_78000_M2 0.050
r 24000_80000_M1 24000_80000_M2 0.050
r 24000_82000_M1 24000_82000_M2 0.050
r 24000_84000_M1 24000_84000_M2 0.050
r 24000_86000_M1 24000_86000_M2 0.050
r 24000_88000_M1 24000_88000_M2 0.050
r 24000_90000_M1 24000_90000_M2 0.050
r 24000_92000_M1 24000_92000_M2 0.050
r 24000_94000_M1 24000_94000_M2 0.050
r 24000_96000_M1 24000_96000_M2 0.050
r 24000_98000_M1 24000_98000_M2 0.050
r 24000_100000_M1 24000_100000_M2 0.050
r 26000_2000_M1 26000_2000_M2 0.050
r 26000_4000_M1 26000_4000_M2 0.050
r 26000_6000_M1 26000_6000_M2 0.050
r 26000_8000_M1 26000_8000_M2 0.050
r 26000_10000_M1 26000_10000_M2 0.050
r 26000_12000_M1 26000_12000_M2 0.050
r 26000_14000_M1 26000_14000_M2 0.050
r 26000_16000_M1 26000_16000_M2 0.050
r 26000_18000_M1 26000_18000_M2 0.050
r 26000_20000_M1 26000_20000_M2 0.050
r 26000_22000_M1 26000_22000_M2 0.050
r 26000_24000_M1 26000_24000_M2 0.050
r 26000_26000_M1 26000_26000_M2 0.050
r 26000_28000_M1 26000_28000_M2 0.050
r 26000_30000_M1 26000_30000_M2 0.050
r 26000_32000_M1 26000_32000_M2 0.050
r 26000_34000_M1 26000_34000_M2 0.050
r 26000_36000_M1 26000_36000_M2 0.050
r 26000_38000_M1 26000_38000_M2 0.050
r 26000_40000_M1 26000_40000_M2 0.050
r 26000_42000_M1 26000_42000_M2 0.050
r 26000_44000_M1 26000_44000_M2 0.050
r 26000_46000_M1 26000_46000_M2 0.050
r 26000_48000_M1 26000_48000_M2 0.050
r 26000_50000_M1 26000_50000_M2 0.050
r 26000_52000_M1 26000_52000_M2 0.050
r 26000_54000_M1 26000_54000_M2 0.050
r 26000_56000_M1 26000_56000_M2 0.050
r 26000_58000_M1 26000_58000_M2 0.050
r 26000_60000_M1 26000_60000_M2 0.050
r 26000_62000_M1 26000_62000_M2 0.050
r 26000_64000_M1 26000_64000_M2 0.050
r 26000_66000_M1 26000_66000_M2 0.050
r 26000_68000_M1 26000_68000_M2 0.050
r 26000_70000_M1 26000_70000_M2 0.050
r 26000_72000_M1 26000_72000_M2 0.050
r 26000_74000_M1 26000_74000_M2 0.050
r 26000_76000_M1 26000_76000_M2 0.050
r 26000_78000_M1 26000_78000_M2 0.050
r 26000_80000_M1 26000_80000_M2 0.050
r 26000_82000_M1 26000_82000_M2 0.050
r 26000_84000_M1 26000_84000_M2 0.050
r 26000_86000_M1 26000_86000_M2 0.050
r 26000_88000_M1 26000_88000_M2 0.050
r 26000_90000_M1 26000_90000_M2 0.050
r 26000_92000_M1 26000_92000_M2 0.050
r 26000_94000_M1 26000_94000_M2 0.050
r 26000_96000_M1 26000_96000_M2 0.050
r 26000_98000_M1 26000_98000_M2 0.050
r 26000_100000_M1 26000_100000_M2 0.050
r 28000_2000_M1 28000_2000_M2 0.050
r 28000_4000_M1 28000_4000_M2 0.050
r 28000_6000_M1 28000_6000_M2 0.050
r 28000_8000_M1 28000_8000_M2 0.050
r 28000_10000_M1 28000_10000_M2 0.050
r 28000_12000_M1 28000_12000_M2 0.050
r 28000_14000_M1 28000_14000_M2 0.050
r 28000_16000_M1 28000_16000_M2 0.050
r 28000_18000_M1 28000_18000_M2 0.050
r 28000_20000_M1 28000_20000_M2 0.050
r 28000_22000_M1 28000_22000_M2 0.050
r 28000_24000_M1 28000_24000_M2 0.050
r 28000_26000_M1 28000_26000_M2 0.050
r 28000_28000_M1 28000_28000_M2 0.050
r 28000_30000_M1 28000_30000_M2 0.050
r 28000_32000_M1 28000_32000_M2 0.050
r 28000_34000_M1 28000_34000_M2 0.050
r 28000_36000_M1 28000_36000_M2 0.050
r 28000_38000_M1 28000_38000_M2 0.050
r 28000_40000_M1 28000_40000_M2 0.050
r 28000_42000_M1 28000_42000_M2 0.050
r 28000_44000_M1 28000_44000_M2 0.050
r 28000_46000_M1 28000_46000_M2 0.050
r 28000_48000_M1 28000_48000_M2 0.050
r 28000_50000_M1 28000_50000_M2 0.050
r 28000_52000_M1 28000_52000_M2 0.050
r 28000_54000_M1 28000_54000_M2 0.050
r 28000_56000_M1 28000_56000_M2 0.050
r 28000_58000_M1 28000_58000_M2 0.050
r 28000_60000_M1 28000_60000_M2 0.050
r 28000_62000_M1 28000_62000_M2 0.050
r 28000_64000_M1 28000_64000_M2 0.050
r 28000_66000_M1 28000_66000_M2 0.050
r 28000_68000_M1 28000_68000_M2 0.050
r 28000_70000_M1 28000_70000_M2 0.050
r 28000_72000_M1 28000_72000_M2 0.050
r 28000_74000_M1 28000_74000_M2 0.050
r 28000_76000_M1 28000_76000_M2 0.050
r 28000_78000_M1 28000_78000_M2 0.050
r 28000_80000_M1 28000_80000_M2 0.050
r 28000_82000_M1 28000_82000_M2 0.050
r 28000_84000_M1 28000_84000_M2 0.050
r 28000_86000_M1 28000_86000_M2 0.050
r 28000_88000_M1 28000_88000_M2 0.050
r 28000_90000_M1 28000_90000_M2 0.050
r 28000_92000_M1 28000_92000_M2 0.050
r 28000_94000_M1 28000_94000_M2 0.050
r 28000_96000_M1 28000_96000_M2 0.050
r 28000_98000_M1 28000_98000_M2 0.050
r 28000_100000_M1 28000_100000_M2 0.050
r 30000_2000_M1 30000_2000_M2 0.050
r 30000_4000_M1 30000_4000_M2 0.050
r 30000_6000_M1 30000_6000_M2 0.050
r 30000_8000_M1 30000_8000_M2 0.050
r 30000_10000_M1 30000_10000_M2 0.050
r 30000_12000_M1 30000_12000_M2 0.050
r 30000_14000_M1 30000_14000_M2 0.050
r 30000_16000_M1 30000_16000_M2 0.050
r 30000_18000_M1 30000_18000_M2 0.050
r 30000_20000_M1 30000_20000_M2 0.050
r 30000_22000_M1 30000_22000_M2 0.050
r 30000_24000_M1 30000_24000_M2 0.050
r 30000_26000_M1 30000_26000_M2 0.050
r 30000_28000_M1 30000_28000_M2 0.050
r 30000_30000_M1 30000_30000_M2 0.050
r 30000_32000_M1 30000_32000_M2 0.050
r 30000_34000_M1 30000_34000_M2 0.050
r 30000_36000_M1 30000_36000_M2 0.050
r 30000_38000_M1 30000_38000_M2 0.050
r 30000_40000_M1 30000_40000_M2 0.050
r 30000_42000_M1 30000_42000_M2 0.050
r 30000_44000_M1 30000_44000_M2 0.050
r 30000_46000_M1 30000_46000_M2 0.050
r 30000_48000_M1 30000_48000_M2 0.050
r 30000_50000_M1 30000_50000_M2 0.050
r 30000_52000_M1 30000_52000_M2 0.050
r 30000_54000_M1 30000_54000_M2 0.050
r 30000_56000_M1 30000_56000_M2 0.050
r 30000_58000_M1 30000_58000_M2 0.050
r 30000_60000_M1 30000_60000_M2 0.050
r 30000_62000_M1 30000_62000_M2 0.050
r 30000_64000_M1 30000_64000_M2 0.050
r 30000_66000_M1 30000_66000_M2 0.050
r 30000_68000_M1 30000_68000_M2 0.050
r 30000_70000_M1 30000_70000_M2 0.050
r 30000_72000_M1 30000_72000_M2 0.050
r 30000_74000_M1 30000_74000_M2 0.050
r 30000_76000_M1 30000_76000_M2 0.050
r 30000_78000_M1 30000_78000_M2 0.050
r 30000_80000_M1 30000_80000_M2 0.050
r 30000_82000_M1 30000_82000_M2 0.050
r 30000_84000_M1 30000_84000_M2 0.050
r 30000_86000_M1 30000_86000_M2 0.050
r 30000_88000_M1 30000_88000_M2 0.050
r 30000_90000_M1 30000_90000_M2 0.050
r 30000_92000_M1 30000_92000_M2 0.050
r 30000_94000_M1 30000_94000_M2 0.050
r 30000_96000_M1 30000_96000_M2 0.050
r 30000_98000_M1 30000_98000_M2 0.050
r 30000_100000_M1 30000_100000_M2 0.050
r 32000_2000_M1 32000_2000_M2 0.050
r 32000_4000_M1 32000_4000_M2 0.050
r 32000_6000_M1 32000_6000_M2 0.050
r 32000_8000_M1 32000_8000_M2 0.050
r 32000_10000_M1 32000_10000_M2 0.050
r 32000_12000_M1 32000_12000_M2 0.050
r 32000_14000_M1 32000_14000_M2 0.050
r 32000_16000_M1 32000_16000_M2 0.050
r 32000_18000_M1 32000_18000_M2 0.050
r 32000_20000_M1 32000_20000_M2 0.050
r 32000_22000_M1 32000_22000_M2 0.050
r 32000_24000_M1 32000_24000_M2 0.050
r 32000_26000_M1 32000_26000_M2 0.050
r 32000_28000_M1 32000_28000_M2 0.050
r 32000_30000_M1 32000_30000_M2 0.050
r 32000_32000_M1 32000_32000_M2 0.050
r 32000_34000_M1 32000_34000_M2 0.050
r 32000_36000_M1 32000_36000_M2 0.050
r 32000_38000_M1 32000_38000_M2 0.050
r 32000_40000_M1 32000_40000_M2 0.050
r 32000_42000_M1 32000_42000_M2 0.050
r 32000_44000_M1 32000_44000_M2 0.050
r 32000_46000_M1 32000_46000_M2 0.050
r 32000_48000_M1 32000_48000_M2 0.050
r 32000_50000_M1 32000_50000_M2 0.050
r 32000_52000_M1 32000_52000_M2 0.050
r 32000_54000_M1 32000_54000_M2 0.050
r 32000_56000_M1 32000_56000_M2 0.050
r 32000_58000_M1 32000_58000_M2 0.050
r 32000_60000_M1 32000_60000_M2 0.050
r 32000_62000_M1 32000_62000_M2 0.050
r 32000_64000_M1 32000_64000_M2 0.050
r 32000_66000_M1 32000_66000_M2 0.050
r 32000_68000_M1 32000_68000_M2 0.050
r 32000_70000_M1 32000_70000_M2 0.050
r 32000_72000_M1 32000_72000_M2 0.050
r 32000_74000_M1 32000_74000_M2 0.050
r 32000_76000_M1 32000_76000_M2 0.050
r 32000_78000_M1 32000_78000_M2 0.050
r 32000_80000_M1 32000_80000_M2 0.050
r 32000_82000_M1 32000_82000_M2 0.050
r 32000_84000_M1 32000_84000_M2 0.050
r 32000_86000_M1 32000_86000_M2 0.050
r 32000_88000_M1 32000_88000_M2 0.050
r 32000_90000_M1 32000_90000_M2 0.050
r 32000_92000_M1 32000_92000_M2 0.050
r 32000_94000_M1 32000_94000_M2 0.050
r 32000_96000_M1 32000_96000_M2 0.050
r 32000_98000_M1 32000_98000_M2 0.050
r 32000_100000_M1 32000_100000_M2 0.050
r 34000_2000_M1 34000_2000_M2 0.050
r 34000_4000_M1 34000_4000_M2 0.050
r 34000_6000_M1 34000_6000_M2 0.050
r 34000_8000_M1 34000_8000_M2 0.050
r 34000_10000_M1 34000_10000_M2 0.050
r 34000_12000_M1 34000_12000_M2 0.050
r 34000_14000_M1 34000_14000_M2 0.050
r 34000_16000_M1 34000_16000_M2 0.050
r 34000_18000_M1 34000_18000_M2 0.050
r 34000_20000_M1 34000_20000_M2 0.050
r 34000_22000_M1 34000_22000_M2 0.050
r 34000_24000_M1 34000_24000_M2 0.050
r 34000_26000_M1 34000_26000_M2 0.050
r 34000_28000_M1 34000_28000_M2 0.050
r 34000_30000_M1 34000_30000_M2 0.050
r 34000_32000_M1 34000_32000_M2 0.050
r 34000_34000_M1 34000_34000_M2 0.050
r 34000_36000_M1 34000_36000_M2 0.050
r 34000_38000_M1 34000_38000_M2 0.050
r 34000_40000_M1 34000_40000_M2 0.050
r 34000_42000_M1 34000_42000_M2 0.050
r 34000_44000_M1 34000_44000_M2 0.050
r 34000_46000_M1 34000_46000_M2 0.050
r 34000_48000_M1 34000_48000_M2 0.050
r 34000_50000_M1 34000_50000_M2 0.050
r 34000_52000_M1 34000_52000_M2 0.050
r 34000_54000_M1 34000_54000_M2 0.050
r 34000_56000_M1 34000_56000_M2 0.050
r 34000_58000_M1 34000_58000_M2 0.050
r 34000_60000_M1 34000_60000_M2 0.050
r 34000_62000_M1 34000_62000_M2 0.050
r 34000_64000_M1 34000_64000_M2 0.050
r 34000_66000_M1 34000_66000_M2 0.050
r 34000_68000_M1 34000_68000_M2 0.050
r 34000_70000_M1 34000_70000_M2 0.050
r 34000_72000_M1 34000_72000_M2 0.050
r 34000_74000_M1 34000_74000_M2 0.050
r 34000_76000_M1 34000_76000_M2 0.050
r 34000_78000_M1 34000_78000_M2 0.050
r 34000_80000_M1 34000_80000_M2 0.050
r 34000_82000_M1 34000_82000_M2 0.050
r 34000_84000_M1 34000_84000_M2 0.050
r 34000_86000_M1 34000_86000_M2 0.050
r 34000_88000_M1 34000_88000_M2 0.050
r 34000_90000_M1 34000_90000_M2 0.050
r 34000_92000_M1 34000_92000_M2 0.050
r 34000_94000_M1 34000_94000_M2 0.050
r 34000_96000_M1 34000_96000_M2 0.050
r 34000_98000_M1 34000_98000_M2 0.050
r 34000_100000_M1 34000_100000_M2 0.050
r 36000_2000_M1 36000_2000_M2 0.050
r 36000_4000_M1 36000_4000_M2 0.050
r 36000_6000_M1 36000_6000_M2 0.050
r 36000_8000_M1 36000_8000_M2 0.050
r 36000_10000_M1 36000_10000_M2 0.050
r 36000_12000_M1 36000_12000_M2 0.050
r 36000_14000_M1 36000_14000_M2 0.050
r 36000_16000_M1 36000_16000_M2 0.050
r 36000_18000_M1 36000_18000_M2 0.050
r 36000_20000_M1 36000_20000_M2 0.050
r 36000_22000_M1 36000_22000_M2 0.050
r 36000_24000_M1 36000_24000_M2 0.050
r 36000_26000_M1 36000_26000_M2 0.050
r 36000_28000_M1 36000_28000_M2 0.050
r 36000_30000_M1 36000_30000_M2 0.050
r 36000_32000_M1 36000_32000_M2 0.050
r 36000_34000_M1 36000_34000_M2 0.050
r 36000_36000_M1 36000_36000_M2 0.050
r 36000_38000_M1 36000_38000_M2 0.050
r 36000_40000_M1 36000_40000_M2 0.050
r 36000_42000_M1 36000_42000_M2 0.050
r 36000_44000_M1 36000_44000_M2 0.050
r 36000_46000_M1 36000_46000_M2 0.050
r 36000_48000_M1 36000_48000_M2 0.050
r 36000_50000_M1 36000_50000_M2 0.050
r 36000_52000_M1 36000_52000_M2 0.050
r 36000_54000_M1 36000_54000_M2 0.050
r 36000_56000_M1 36000_56000_M2 0.050
r 36000_58000_M1 36000_58000_M2 0.050
r 36000_60000_M1 36000_60000_M2 0.050
r 36000_62000_M1 36000_62000_M2 0.050
r 36000_64000_M1 36000_64000_M2 0.050
r 36000_66000_M1 36000_66000_M2 0.050
r 36000_68000_M1 36000_68000_M2 0.050
r 36000_70000_M1 36000_70000_M2 0.050
r 36000_72000_M1 36000_72000_M2 0.050
r 36000_74000_M1 36000_74000_M2 0.050
r 36000_76000_M1 36000_76000_M2 0.050
r 36000_78000_M1 36000_78000_M2 0.050
r 36000_80000_M1 36000_80000_M2 0.050
r 36000_82000_M1 36000_82000_M2 0.050
r 36000_84000_M1 36000_84000_M2 0.050
r 36000_86000_M1 36000_86000_M2 0.050
r 36000_88000_M1 36000_88000_M2 0.050
r 36000_90000_M1 36000_90000_M2 0.050
r 36000_92000_M1 36000_92000_M2 0.050
r 36000_94000_M1 36000_94000_M2 0.050
r 36000_96000_M1 36000_96000_M2 0.050
r 36000_98000_M1 36000_98000_M2 0.050
r 36000_100000_M1 36000_100000_M2 0.050
r 38000_2000_M1 38000_2000_M2 0.050
r 38000_4000_M1 38000_4000_M2 0.050
r 38000_6000_M1 38000_6000_M2 0.050
r 38000_8000_M1 38000_8000_M2 0.050
r 38000_10000_M1 38000_10000_M2 0.050
r 38000_12000_M1 38000_12000_M2 0.050
r 38000_14000_M1 38000_14000_M2 0.050
r 38000_16000_M1 38000_16000_M2 0.050
r 38000_18000_M1 38000_18000_M2 0.050
r 38000_20000_M1 38000_20000_M2 0.050
r 38000_22000_M1 38000_22000_M2 0.050
r 38000_24000_M1 38000_24000_M2 0.050
r 38000_26000_M1 38000_26000_M2 0.050
r 38000_28000_M1 38000_28000_M2 0.050
r 38000_30000_M1 38000_30000_M2 0.050
r 38000_32000_M1 38000_32000_M2 0.050
r 38000_34000_M1 38000_34000_M2 0.050
r 38000_36000_M1 38000_36000_M2 0.050
r 38000_38000_M1 38000_38000_M2 0.050
r 38000_40000_M1 38000_40000_M2 0.050
r 38000_42000_M1 38000_42000_M2 0.050
r 38000_44000_M1 38000_44000_M2 0.050
r 38000_46000_M1 38000_46000_M2 0.050
r 38000_48000_M1 38000_48000_M2 0.050
r 38000_50000_M1 38000_50000_M2 0.050
r 38000_52000_M1 38000_52000_M2 0.050
r 38000_54000_M1 38000_54000_M2 0.050
r 38000_56000_M1 38000_56000_M2 0.050
r 38000_58000_M1 38000_58000_M2 0.050
r 38000_60000_M1 38000_60000_M2 0.050
r 38000_62000_M1 38000_62000_M2 0.050
r 38000_64000_M1 38000_64000_M2 0.050
r 38000_66000_M1 38000_66000_M2 0.050
r 38000_68000_M1 38000_68000_M2 0.050
r 38000_70000_M1 38000_70000_M2 0.050
r 38000_72000_M1 38000_72000_M2 0.050
r 38000_74000_M1 38000_74000_M2 0.050
r 38000_76000_M1 38000_76000_M2 0.050
r 38000_78000_M1 38000_78000_M2 0.050
r 38000_80000_M1 38000_80000_M2 0.050
r 38000_82000_M1 38000_82000_M2 0.050
r 38000_84000_M1 38000_84000_M2 0.050
r 38000_86000_M1 38000_86000_M2 0.050
r 38000_88000_M1 38000_88000_M2 0.050
r 38000_90000_M1 38000_90000_M2 0.050
r 38000_92000_M1 38000_92000_M2 0.050
r 38000_94000_M1 38000_94000_M2 0.050
r 38000_96000_M1 38000_96000_M2 0.050
r 38000_98000_M1 38000_98000_M2 0.050
r 38000_100000_M1 38000_100000_M2 0.050
r 40000_2000_M1 40000_2000_M2 0.050
r 40000_4000_M1 40000_4000_M2 0.050
r 40000_6000_M1 40000_6000_M2 0.050
r 40000_8000_M1 40000_8000_M2 0.050
r 40000_10000_M1 40000_10000_M2 0.050
r 40000_12000_M1 40000_12000_M2 0.050
r 40000_14000_M1 40000_14000_M2 0.050
r 40000_16000_M1 40000_16000_M2 0.050
r 40000_18000_M1 40000_18000_M2 0.050
r 40000_20000_M1 40000_20000_M2 0.050
r 40000_22000_M1 40000_22000_M2 0.050
r 40000_24000_M1 40000_24000_M2 0.050
r 40000_26000_M1 40000_26000_M2 0.050
r 40000_28000_M1 40000_28000_M2 0.050
r 40000_30000_M1 40000_30000_M2 0.050
r 40000_32000_M1 40000_32000_M2 0.050
r 40000_34000_M1 40000_34000_M2 0.050
r 40000_36000_M1 40000_36000_M2 0.050
r 40000_38000_M1 40000_38000_M2 0.050
r 40000_40000_M1 40000_40000_M2 0.050
r 40000_42000_M1 40000_42000_M2 0.050
r 40000_44000_M1 40000_44000_M2 0.050
r 40000_46000_M1 40000_46000_M2 0.050
r 40000_48000_M1 40000_48000_M2 0.050
r 40000_50000_M1 40000_50000_M2 0.050
r 40000_52000_M1 40000_52000_M2 0.050
r 40000_54000_M1 40000_54000_M2 0.050
r 40000_56000_M1 40000_56000_M2 0.050
r 40000_58000_M1 40000_58000_M2 0.050
r 40000_60000_M1 40000_60000_M2 0.050
r 40000_62000_M1 40000_62000_M2 0.050
r 40000_64000_M1 40000_64000_M2 0.050
r 40000_66000_M1 40000_66000_M2 0.050
r 40000_68000_M1 40000_68000_M2 0.050
r 40000_70000_M1 40000_70000_M2 0.050
r 40000_72000_M1 40000_72000_M2 0.050
r 40000_74000_M1 40000_74000_M2 0.050
r 40000_76000_M1 40000_76000_M2 0.050
r 40000_78000_M1 40000_78000_M2 0.050
r 40000_80000_M1 40000_80000_M2 0.050
r 40000_82000_M1 40000_82000_M2 0.050
r 40000_84000_M1 40000_84000_M2 0.050
r 40000_86000_M1 40000_86000_M2 0.050
r 40000_88000_M1 40000_88000_M2 0.050
r 40000_90000_M1 40000_90000_M2 0.050
r 40000_92000_M1 40000_92000_M2 0.050
r 40000_94000_M1 40000_94000_M2 0.050
r 40000_96000_M1 40000_96000_M2 0.050
r 40000_98000_M1 40000_98000_M2 0.050
r 40000_100000_M1 40000_100000_M2 0.050
r 42000_2000_M1 42000_2000_M2 0.050
r 42000_4000_M1 42000_4000_M2 0.050
r 42000_6000_M1 42000_6000_M2 0.050
r 42000_8000_M1 42000_8000_M2 0.050
r 42000_10000_M1 42000_10000_M2 0.050
r 42000_12000_M1 42000_12000_M2 0.050
r 42000_14000_M1 42000_14000_M2 0.050
r 42000_16000_M1 42000_16000_M2 0.050
r 42000_18000_M1 42000_18000_M2 0.050
r 42000_20000_M1 42000_20000_M2 0.050
r 42000_22000_M1 42000_22000_M2 0.050
r 42000_24000_M1 42000_24000_M2 0.050
r 42000_26000_M1 42000_26000_M2 0.050
r 42000_28000_M1 42000_28000_M2 0.050
r 42000_30000_M1 42000_30000_M2 0.050
r 42000_32000_M1 42000_32000_M2 0.050
r 42000_34000_M1 42000_34000_M2 0.050
r 42000_36000_M1 42000_36000_M2 0.050
r 42000_38000_M1 42000_38000_M2 0.050
r 42000_40000_M1 42000_40000_M2 0.050
r 42000_42000_M1 42000_42000_M2 0.050
r 42000_44000_M1 42000_44000_M2 0.050
r 42000_46000_M1 42000_46000_M2 0.050
r 42000_48000_M1 42000_48000_M2 0.050
r 42000_50000_M1 42000_50000_M2 0.050
r 42000_52000_M1 42000_52000_M2 0.050
r 42000_54000_M1 42000_54000_M2 0.050
r 42000_56000_M1 42000_56000_M2 0.050
r 42000_58000_M1 42000_58000_M2 0.050
r 42000_60000_M1 42000_60000_M2 0.050
r 42000_62000_M1 42000_62000_M2 0.050
r 42000_64000_M1 42000_64000_M2 0.050
r 42000_66000_M1 42000_66000_M2 0.050
r 42000_68000_M1 42000_68000_M2 0.050
r 42000_70000_M1 42000_70000_M2 0.050
r 42000_72000_M1 42000_72000_M2 0.050
r 42000_74000_M1 42000_74000_M2 0.050
r 42000_76000_M1 42000_76000_M2 0.050
r 42000_78000_M1 42000_78000_M2 0.050
r 42000_80000_M1 42000_80000_M2 0.050
r 42000_82000_M1 42000_82000_M2 0.050
r 42000_84000_M1 42000_84000_M2 0.050
r 42000_86000_M1 42000_86000_M2 0.050
r 42000_88000_M1 42000_88000_M2 0.050
r 42000_90000_M1 42000_90000_M2 0.050
r 42000_92000_M1 42000_92000_M2 0.050
r 42000_94000_M1 42000_94000_M2 0.050
r 42000_96000_M1 42000_96000_M2 0.050
r 42000_98000_M1 42000_98000_M2 0.050
r 42000_100000_M1 42000_100000_M2 0.050
r 44000_2000_M1 44000_2000_M2 0.050
r 44000_4000_M1 44000_4000_M2 0.050
r 44000_6000_M1 44000_6000_M2 0.050
r 44000_8000_M1 44000_8000_M2 0.050
r 44000_10000_M1 44000_10000_M2 0.050
r 44000_12000_M1 44000_12000_M2 0.050
r 44000_14000_M1 44000_14000_M2 0.050
r 44000_16000_M1 44000_16000_M2 0.050
r 44000_18000_M1 44000_18000_M2 0.050
r 44000_20000_M1 44000_20000_M2 0.050
r 44000_22000_M1 44000_22000_M2 0.050
r 44000_24000_M1 44000_24000_M2 0.050
r 44000_26000_M1 44000_26000_M2 0.050
r 44000_28000_M1 44000_28000_M2 0.050
r 44000_30000_M1 44000_30000_M2 0.050
r 44000_32000_M1 44000_32000_M2 0.050
r 44000_34000_M1 44000_34000_M2 0.050
r 44000_36000_M1 44000_36000_M2 0.050
r 44000_38000_M1 44000_38000_M2 0.050
r 44000_40000_M1 44000_40000_M2 0.050
r 44000_42000_M1 44000_42000_M2 0.050
r 44000_44000_M1 44000_44000_M2 0.050
r 44000_46000_M1 44000_46000_M2 0.050
r 44000_48000_M1 44000_48000_M2 0.050
r 44000_50000_M1 44000_50000_M2 0.050
r 44000_52000_M1 44000_52000_M2 0.050
r 44000_54000_M1 44000_54000_M2 0.050
r 44000_56000_M1 44000_56000_M2 0.050
r 44000_58000_M1 44000_58000_M2 0.050
r 44000_60000_M1 44000_60000_M2 0.050
r 44000_62000_M1 44000_62000_M2 0.050
r 44000_64000_M1 44000_64000_M2 0.050
r 44000_66000_M1 44000_66000_M2 0.050
r 44000_68000_M1 44000_68000_M2 0.050
r 44000_70000_M1 44000_70000_M2 0.050
r 44000_72000_M1 44000_72000_M2 0.050
r 44000_74000_M1 44000_74000_M2 0.050
r 44000_76000_M1 44000_76000_M2 0.050
r 44000_78000_M1 44000_78000_M2 0.050
r 44000_80000_M1 44000_80000_M2 0.050
r 44000_82000_M1 44000_82000_M2 0.050
r 44000_84000_M1 44000_84000_M2 0.050
r 44000_86000_M1 44000_86000_M2 0.050
r 44000_88000_M1 44000_88000_M2 0.050
r 44000_90000_M1 44000_90000_M2 0.050
r 44000_92000_M1 44000_92000_M2 0.050
r 44000_94000_M1 44000_94000_M2 0.050
r 44000_96000_M1 44000_96000_M2 0.050
r 44000_98000_M1 44000_98000_M2 0.050
r 44000_100000_M1 44000_100000_M2 0.050
r 46000_2000_M1 46000_2000_M2 0.050
r 46000_4000_M1 46000_4000_M2 0.050
r 46000_6000_M1 46000_6000_M2 0.050
r 46000_8000_M1 46000_8000_M2 0.050
r 46000_10000_M1 46000_10000_M2 0.050
r 46000_12000_M1 46000_12000_M2 0.050
r 46000_14000_M1 46000_14000_M2 0.050
r 46000_16000_M1 46000_16000_M2 0.050
r 46000_18000_M1 46000_18000_M2 0.050
r 46000_20000_M1 46000_20000_M2 0.050
r 46000_22000_M1 46000_22000_M2 0.050
r 46000_24000_M1 46000_24000_M2 0.050
r 46000_26000_M1 46000_26000_M2 0.050
r 46000_28000_M1 46000_28000_M2 0.050
r 46000_30000_M1 46000_30000_M2 0.050
r 46000_32000_M1 46000_32000_M2 0.050
r 46000_34000_M1 46000_34000_M2 0.050
r 46000_36000_M1 46000_36000_M2 0.050
r 46000_38000_M1 46000_38000_M2 0.050
r 46000_40000_M1 46000_40000_M2 0.050
r 46000_42000_M1 46000_42000_M2 0.050
r 46000_44000_M1 46000_44000_M2 0.050
r 46000_46000_M1 46000_46000_M2 0.050
r 46000_48000_M1 46000_48000_M2 0.050
r 46000_50000_M1 46000_50000_M2 0.050
r 46000_52000_M1 46000_52000_M2 0.050
r 46000_54000_M1 46000_54000_M2 0.050
r 46000_56000_M1 46000_56000_M2 0.050
r 46000_58000_M1 46000_58000_M2 0.050
r 46000_60000_M1 46000_60000_M2 0.050
r 46000_62000_M1 46000_62000_M2 0.050
r 46000_64000_M1 46000_64000_M2 0.050
r 46000_66000_M1 46000_66000_M2 0.050
r 46000_68000_M1 46000_68000_M2 0.050
r 46000_70000_M1 46000_70000_M2 0.050
r 46000_72000_M1 46000_72000_M2 0.050
r 46000_74000_M1 46000_74000_M2 0.050
r 46000_76000_M1 46000_76000_M2 0.050
r 46000_78000_M1 46000_78000_M2 0.050
r 46000_80000_M1 46000_80000_M2 0.050
r 46000_82000_M1 46000_82000_M2 0.050
r 46000_84000_M1 46000_84000_M2 0.050
r 46000_86000_M1 46000_86000_M2 0.050
r 46000_88000_M1 46000_88000_M2 0.050
r 46000_90000_M1 46000_90000_M2 0.050
r 46000_92000_M1 46000_92000_M2 0.050
r 46000_94000_M1 46000_94000_M2 0.050
r 46000_96000_M1 46000_96000_M2 0.050
r 46000_98000_M1 46000_98000_M2 0.050
r 46000_100000_M1 46000_100000_M2 0.050
r 48000_2000_M1 48000_2000_M2 0.050
r 48000_4000_M1 48000_4000_M2 0.050
r 48000_6000_M1 48000_6000_M2 0.050
r 48000_8000_M1 48000_8000_M2 0.050
r 48000_10000_M1 48000_10000_M2 0.050
r 48000_12000_M1 48000_12000_M2 0.050
r 48000_14000_M1 48000_14000_M2 0.050
r 48000_16000_M1 48000_16000_M2 0.050
r 48000_18000_M1 48000_18000_M2 0.050
r 48000_20000_M1 48000_20000_M2 0.050
r 48000_22000_M1 48000_22000_M2 0.050
r 48000_24000_M1 48000_24000_M2 0.050
r 48000_26000_M1 48000_26000_M2 0.050
r 48000_28000_M1 48000_28000_M2 0.050
r 48000_30000_M1 48000_30000_M2 0.050
r 48000_32000_M1 48000_32000_M2 0.050
r 48000_34000_M1 48000_34000_M2 0.050
r 48000_36000_M1 48000_36000_M2 0.050
r 48000_38000_M1 48000_38000_M2 0.050
r 48000_40000_M1 48000_40000_M2 0.050
r 48000_42000_M1 48000_42000_M2 0.050
r 48000_44000_M1 48000_44000_M2 0.050
r 48000_46000_M1 48000_46000_M2 0.050
r 48000_48000_M1 48000_48000_M2 0.050
r 48000_50000_M1 48000_50000_M2 0.050
r 48000_52000_M1 48000_52000_M2 0.050
r 48000_54000_M1 48000_54000_M2 0.050
r 48000_56000_M1 48000_56000_M2 0.050
r 48000_58000_M1 48000_58000_M2 0.050
r 48000_60000_M1 48000_60000_M2 0.050
r 48000_62000_M1 48000_62000_M2 0.050
r 48000_64000_M1 48000_64000_M2 0.050
r 48000_66000_M1 48000_66000_M2 0.050
r 48000_68000_M1 48000_68000_M2 0.050
r 48000_70000_M1 48000_70000_M2 0.050
r 48000_72000_M1 48000_72000_M2 0.050
r 48000_74000_M1 48000_74000_M2 0.050
r 48000_76000_M1 48000_76000_M2 0.050
r 48000_78000_M1 48000_78000_M2 0.050
r 48000_80000_M1 48000_80000_M2 0.050
r 48000_82000_M1 48000_82000_M2 0.050
r 48000_84000_M1 48000_84000_M2 0.050
r 48000_86000_M1 48000_86000_M2 0.050
r 48000_88000_M1 48000_88000_M2 0.050
r 48000_90000_M1 48000_90000_M2 0.050
r 48000_92000_M1 48000_92000_M2 0.050
r 48000_94000_M1 48000_94000_M2 0.050
r 48000_96000_M1 48000_96000_M2 0.050
r 48000_98000_M1 48000_98000_M2 0.050
r 48000_100000_M1 48000_100000_M2 0.050
r 50000_2000_M1 50000_2000_M2 0.050
r 50000_4000_M1 50000_4000_M2 0.050
r 50000_6000_M1 50000_6000_M2 0.050
r 50000_8000_M1 50000_8000_M2 0.050
r 50000_10000_M1 50000_10000_M2 0.050
r 50000_12000_M1 50000_12000_M2 0.050
r 50000_14000_M1 50000_14000_M2 0.050
r 50000_16000_M1 50000_16000_M2 0.050
r 50000_18000_M1 50000_18000_M2 0.050
r 50000_20000_M1 50000_20000_M2 0.050
r 50000_22000_M1 50000_22000_M2 0.050
r 50000_24000_M1 50000_24000_M2 0.050
r 50000_26000_M1 50000_26000_M2 0.050
r 50000_28000_M1 50000_28000_M2 0.050
r 50000_30000_M1 50000_30000_M2 0.050
r 50000_32000_M1 50000_32000_M2 0.050
r 50000_34000_M1 50000_34000_M2 0.050
r 50000_36000_M1 50000_36000_M2 0.050
r 50000_38000_M1 50000_38000_M2 0.050
r 50000_40000_M1 50000_40000_M2 0.050
r 50000_42000_M1 50000_42000_M2 0.050
r 50000_44000_M1 50000_44000_M2 0.050
r 50000_46000_M1 50000_46000_M2 0.050
r 50000_48000_M1 50000_48000_M2 0.050
r 50000_50000_M1 50000_50000_M2 0.050
r 50000_52000_M1 50000_52000_M2 0.050
r 50000_54000_M1 50000_54000_M2 0.050
r 50000_56000_M1 50000_56000_M2 0.050
r 50000_58000_M1 50000_58000_M2 0.050
r 50000_60000_M1 50000_60000_M2 0.050
r 50000_62000_M1 50000_62000_M2 0.050
r 50000_64000_M1 50000_64000_M2 0.050
r 50000_66000_M1 50000_66000_M2 0.050
r 50000_68000_M1 50000_68000_M2 0.050
r 50000_70000_M1 50000_70000_M2 0.050
r 50000_72000_M1 50000_72000_M2 0.050
r 50000_74000_M1 50000_74000_M2 0.050
r 50000_76000_M1 50000_76000_M2 0.050
r 50000_78000_M1 50000_78000_M2 0.050
r 50000_80000_M1 50000_80000_M2 0.050
r 50000_82000_M1 50000_82000_M2 0.050
r 50000_84000_M1 50000_84000_M2 0.050
r 50000_86000_M1 50000_86000_M2 0.050
r 50000_88000_M1 50000_88000_M2 0.050
r 50000_90000_M1 50000_90000_M2 0.050
r 50000_92000_M1 50000_92000_M2 0.050
r 50000_94000_M1 50000_94000_M2 0.050
r 50000_96000_M1 50000_96000_M2 0.050
r 50000_98000_M1 50000_98000_M2 0.050
r 50000_100000_M1 50000_100000_M2 0.050
r 52000_2000_M1 52000_2000_M2 0.050
r 52000_4000_M1 52000_4000_M2 0.050
r 52000_6000_M1 52000_6000_M2 0.050
r 52000_8000_M1 52000_8000_M2 0.050
r 52000_10000_M1 52000_10000_M2 0.050
r 52000_12000_M1 52000_12000_M2 0.050
r 52000_14000_M1 52000_14000_M2 0.050
r 52000_16000_M1 52000_16000_M2 0.050
r 52000_18000_M1 52000_18000_M2 0.050
r 52000_20000_M1 52000_20000_M2 0.050
r 52000_22000_M1 52000_22000_M2 0.050
r 52000_24000_M1 52000_24000_M2 0.050
r 52000_26000_M1 52000_26000_M2 0.050
r 52000_28000_M1 52000_28000_M2 0.050
r 52000_30000_M1 52000_30000_M2 0.050
r 52000_32000_M1 52000_32000_M2 0.050
r 52000_34000_M1 52000_34000_M2 0.050
r 52000_36000_M1 52000_36000_M2 0.050
r 52000_38000_M1 52000_38000_M2 0.050
r 52000_40000_M1 52000_40000_M2 0.050
r 52000_42000_M1 52000_42000_M2 0.050
r 52000_44000_M1 52000_44000_M2 0.050
r 52000_46000_M1 52000_46000_M2 0.050
r 52000_48000_M1 52000_48000_M2 0.050
r 52000_50000_M1 52000_50000_M2 0.050
r 52000_52000_M1 52000_52000_M2 0.050
r 52000_54000_M1 52000_54000_M2 0.050
r 52000_56000_M1 52000_56000_M2 0.050
r 52000_58000_M1 52000_58000_M2 0.050
r 52000_60000_M1 52000_60000_M2 0.050
r 52000_62000_M1 52000_62000_M2 0.050
r 52000_64000_M1 52000_64000_M2 0.050
r 52000_66000_M1 52000_66000_M2 0.050
r 52000_68000_M1 52000_68000_M2 0.050
r 52000_70000_M1 52000_70000_M2 0.050
r 52000_72000_M1 52000_72000_M2 0.050
r 52000_74000_M1 52000_74000_M2 0.050
r 52000_76000_M1 52000_76000_M2 0.050
r 52000_78000_M1 52000_78000_M2 0.050
r 52000_80000_M1 52000_80000_M2 0.050
r 52000_82000_M1 52000_82000_M2 0.050
r 52000_84000_M1 52000_84000_M2 0.050
r 52000_86000_M1 52000_86000_M2 0.050
r 52000_88000_M1 52000_88000_M2 0.050
r 52000_90000_M1 52000_90000_M2 0.050
r 52000_92000_M1 52000_92000_M2 0.050
r 52000_94000_M1 52000_94000_M2 0.050
r 52000_96000_M1 52000_96000_M2 0.050
r 52000_98000_M1 52000_98000_M2 0.050
r 52000_100000_M1 52000_100000_M2 0.050
r 54000_2000_M1 54000_2000_M2 0.050
r 54000_4000_M1 54000_4000_M2 0.050
r 54000_6000_M1 54000_6000_M2 0.050
r 54000_8000_M1 54000_8000_M2 0.050
r 54000_10000_M1 54000_10000_M2 0.050
r 54000_12000_M1 54000_12000_M2 0.050
r 54000_14000_M1 54000_14000_M2 0.050
r 54000_16000_M1 54000_16000_M2 0.050
r 54000_18000_M1 54000_18000_M2 0.050
r 54000_20000_M1 54000_20000_M2 0.050
r 54000_22000_M1 54000_22000_M2 0.050
r 54000_24000_M1 54000_24000_M2 0.050
r 54000_26000_M1 54000_26000_M2 0.050
r 54000_28000_M1 54000_28000_M2 0.050
r 54000_30000_M1 54000_30000_M2 0.050
r 54000_32000_M1 54000_32000_M2 0.050
r 54000_34000_M1 54000_34000_M2 0.050
r 54000_36000_M1 54000_36000_M2 0.050
r 54000_38000_M1 54000_38000_M2 0.050
r 54000_40000_M1 54000_40000_M2 0.050
r 54000_42000_M1 54000_42000_M2 0.050
r 54000_44000_M1 54000_44000_M2 0.050
r 54000_46000_M1 54000_46000_M2 0.050
r 54000_48000_M1 54000_48000_M2 0.050
r 54000_50000_M1 54000_50000_M2 0.050
r 54000_52000_M1 54000_52000_M2 0.050
r 54000_54000_M1 54000_54000_M2 0.050
r 54000_56000_M1 54000_56000_M2 0.050
r 54000_58000_M1 54000_58000_M2 0.050
r 54000_60000_M1 54000_60000_M2 0.050
r 54000_62000_M1 54000_62000_M2 0.050
r 54000_64000_M1 54000_64000_M2 0.050
r 54000_66000_M1 54000_66000_M2 0.050
r 54000_68000_M1 54000_68000_M2 0.050
r 54000_70000_M1 54000_70000_M2 0.050
r 54000_72000_M1 54000_72000_M2 0.050
r 54000_74000_M1 54000_74000_M2 0.050
r 54000_76000_M1 54000_76000_M2 0.050
r 54000_78000_M1 54000_78000_M2 0.050
r 54000_80000_M1 54000_80000_M2 0.050
r 54000_82000_M1 54000_82000_M2 0.050
r 54000_84000_M1 54000_84000_M2 0.050
r 54000_86000_M1 54000_86000_M2 0.050
r 54000_88000_M1 54000_88000_M2 0.050
r 54000_90000_M1 54000_90000_M2 0.050
r 54000_92000_M1 54000_92000_M2 0.050
r 54000_94000_M1 54000_94000_M2 0.050
r 54000_96000_M1 54000_96000_M2 0.050
r 54000_98000_M1 54000_98000_M2 0.050
r 54000_100000_M1 54000_100000_M2 0.050
r 56000_2000_M1 56000_2000_M2 0.050
r 56000_4000_M1 56000_4000_M2 0.050
r 56000_6000_M1 56000_6000_M2 0.050
r 56000_8000_M1 56000_8000_M2 0.050
r 56000_10000_M1 56000_10000_M2 0.050
r 56000_12000_M1 56000_12000_M2 0.050
r 56000_14000_M1 56000_14000_M2 0.050
r 56000_16000_M1 56000_16000_M2 0.050
r 56000_18000_M1 56000_18000_M2 0.050
r 56000_20000_M1 56000_20000_M2 0.050
r 56000_22000_M1 56000_22000_M2 0.050
r 56000_24000_M1 56000_24000_M2 0.050
r 56000_26000_M1 56000_26000_M2 0.050
r 56000_28000_M1 56000_28000_M2 0.050
r 56000_30000_M1 56000_30000_M2 0.050
r 56000_32000_M1 56000_32000_M2 0.050
r 56000_34000_M1 56000_34000_M2 0.050
r 56000_36000_M1 56000_36000_M2 0.050
r 56000_38000_M1 56000_38000_M2 0.050
r 56000_40000_M1 56000_40000_M2 0.050
r 56000_42000_M1 56000_42000_M2 0.050
r 56000_44000_M1 56000_44000_M2 0.050
r 56000_46000_M1 56000_46000_M2 0.050
r 56000_48000_M1 56000_48000_M2 0.050
r 56000_50000_M1 56000_50000_M2 0.050
r 56000_52000_M1 56000_52000_M2 0.050
r 56000_54000_M1 56000_54000_M2 0.050
r 56000_56000_M1 56000_56000_M2 0.050
r 56000_58000_M1 56000_58000_M2 0.050
r 56000_60000_M1 56000_60000_M2 0.050
r 56000_62000_M1 56000_62000_M2 0.050
r 56000_64000_M1 56000_64000_M2 0.050
r 56000_66000_M1 56000_66000_M2 0.050
r 56000_68000_M1 56000_68000_M2 0.050
r 56000_70000_M1 56000_70000_M2 0.050
r 56000_72000_M1 56000_72000_M2 0.050
r 56000_74000_M1 56000_74000_M2 0.050
r 56000_76000_M1 56000_76000_M2 0.050
r 56000_78000_M1 56000_78000_M2 0.050
r 56000_80000_M1 56000_80000_M2 0.050
r 56000_82000_M1 56000_82000_M2 0.050
r 56000_84000_M1 56000_84000_M2 0.050
r 56000_86000_M1 56000_86000_M2 0.050
r 56000_88000_M1 56000_88000_M2 0.050
r 56000_90000_M1 56000_90000_M2 0.050
r 56000_92000_M1 56000_92000_M2 0.050
r 56000_94000_M1 56000_94000_M2 0.050
r 56000_96000_M1 56000_96000_M2 0.050
r 56000_98000_M1 56000_98000_M2 0.050
r 56000_100000_M1 56000_100000_M2 0.050
r 58000_2000_M1 58000_2000_M2 0.050
r 58000_4000_M1 58000_4000_M2 0.050
r 58000_6000_M1 58000_6000_M2 0.050
r 58000_8000_M1 58000_8000_M2 0.050
r 58000_10000_M1 58000_10000_M2 0.050
r 58000_12000_M1 58000_12000_M2 0.050
r 58000_14000_M1 58000_14000_M2 0.050
r 58000_16000_M1 58000_16000_M2 0.050
r 58000_18000_M1 58000_18000_M2 0.050
r 58000_20000_M1 58000_20000_M2 0.050
r 58000_22000_M1 58000_22000_M2 0.050
r 58000_24000_M1 58000_24000_M2 0.050
r 58000_26000_M1 58000_26000_M2 0.050
r 58000_28000_M1 58000_28000_M2 0.050
r 58000_30000_M1 58000_30000_M2 0.050
r 58000_32000_M1 58000_32000_M2 0.050
r 58000_34000_M1 58000_34000_M2 0.050
r 58000_36000_M1 58000_36000_M2 0.050
r 58000_38000_M1 58000_38000_M2 0.050
r 58000_40000_M1 58000_40000_M2 0.050
r 58000_42000_M1 58000_42000_M2 0.050
r 58000_44000_M1 58000_44000_M2 0.050
r 58000_46000_M1 58000_46000_M2 0.050
r 58000_48000_M1 58000_48000_M2 0.050
r 58000_50000_M1 58000_50000_M2 0.050
r 58000_52000_M1 58000_52000_M2 0.050
r 58000_54000_M1 58000_54000_M2 0.050
r 58000_56000_M1 58000_56000_M2 0.050
r 58000_58000_M1 58000_58000_M2 0.050
r 58000_60000_M1 58000_60000_M2 0.050
r 58000_62000_M1 58000_62000_M2 0.050
r 58000_64000_M1 58000_64000_M2 0.050
r 58000_66000_M1 58000_66000_M2 0.050
r 58000_68000_M1 58000_68000_M2 0.050
r 58000_70000_M1 58000_70000_M2 0.050
r 58000_72000_M1 58000_72000_M2 0.050
r 58000_74000_M1 58000_74000_M2 0.050
r 58000_76000_M1 58000_76000_M2 0.050
r 58000_78000_M1 58000_78000_M2 0.050
r 58000_80000_M1 58000_80000_M2 0.050
r 58000_82000_M1 58000_82000_M2 0.050
r 58000_84000_M1 58000_84000_M2 0.050
r 58000_86000_M1 58000_86000_M2 0.050
r 58000_88000_M1 58000_88000_M2 0.050
r 58000_90000_M1 58000_90000_M2 0.050
r 58000_92000_M1 58000_92000_M2 0.050
r 58000_94000_M1 58000_94000_M2 0.050
r 58000_96000_M1 58000_96000_M2 0.050
r 58000_98000_M1 58000_98000_M2 0.050
r 58000_100000_M1 58000_100000_M2 0.050
r 60000_2000_M1 60000_2000_M2 0.050
r 60000_4000_M1 60000_4000_M2 0.050
r 60000_6000_M1 60000_6000_M2 0.050
r 60000_8000_M1 60000_8000_M2 0.050
r 60000_10000_M1 60000_10000_M2 0.050
r 60000_12000_M1 60000_12000_M2 0.050
r 60000_14000_M1 60000_14000_M2 0.050
r 60000_16000_M1 60000_16000_M2 0.050
r 60000_18000_M1 60000_18000_M2 0.050
r 60000_20000_M1 60000_20000_M2 0.050
r 60000_22000_M1 60000_22000_M2 0.050
r 60000_24000_M1 60000_24000_M2 0.050
r 60000_26000_M1 60000_26000_M2 0.050
r 60000_28000_M1 60000_28000_M2 0.050
r 60000_30000_M1 60000_30000_M2 0.050
r 60000_32000_M1 60000_32000_M2 0.050
r 60000_34000_M1 60000_34000_M2 0.050
r 60000_36000_M1 60000_36000_M2 0.050
r 60000_38000_M1 60000_38000_M2 0.050
r 60000_40000_M1 60000_40000_M2 0.050
r 60000_42000_M1 60000_42000_M2 0.050
r 60000_44000_M1 60000_44000_M2 0.050
r 60000_46000_M1 60000_46000_M2 0.050
r 60000_48000_M1 60000_48000_M2 0.050
r 60000_50000_M1 60000_50000_M2 0.050
r 60000_52000_M1 60000_52000_M2 0.050
r 60000_54000_M1 60000_54000_M2 0.050
r 60000_56000_M1 60000_56000_M2 0.050
r 60000_58000_M1 60000_58000_M2 0.050
r 60000_60000_M1 60000_60000_M2 0.050
r 60000_62000_M1 60000_62000_M2 0.050
r 60000_64000_M1 60000_64000_M2 0.050
r 60000_66000_M1 60000_66000_M2 0.050
r 60000_68000_M1 60000_68000_M2 0.050
r 60000_70000_M1 60000_70000_M2 0.050
r 60000_72000_M1 60000_72000_M2 0.050
r 60000_74000_M1 60000_74000_M2 0.050
r 60000_76000_M1 60000_76000_M2 0.050
r 60000_78000_M1 60000_78000_M2 0.050
r 60000_80000_M1 60000_80000_M2 0.050
r 60000_82000_M1 60000_82000_M2 0.050
r 60000_84000_M1 60000_84000_M2 0.050
r 60000_86000_M1 60000_86000_M2 0.050
r 60000_88000_M1 60000_88000_M2 0.050
r 60000_90000_M1 60000_90000_M2 0.050
r 60000_92000_M1 60000_92000_M2 0.050
r 60000_94000_M1 60000_94000_M2 0.050
r 60000_96000_M1 60000_96000_M2 0.050
r 60000_98000_M1 60000_98000_M2 0.050
r 60000_100000_M1 60000_100000_M2 0.050
r 62000_2000_M1 62000_2000_M2 0.050
r 62000_4000_M1 62000_4000_M2 0.050
r 62000_6000_M1 62000_6000_M2 0.050
r 62000_8000_M1 62000_8000_M2 0.050
r 62000_10000_M1 62000_10000_M2 0.050
r 62000_12000_M1 62000_12000_M2 0.050
r 62000_14000_M1 62000_14000_M2 0.050
r 62000_16000_M1 62000_16000_M2 0.050
r 62000_18000_M1 62000_18000_M2 0.050
r 62000_20000_M1 62000_20000_M2 0.050
r 62000_22000_M1 62000_22000_M2 0.050
r 62000_24000_M1 62000_24000_M2 0.050
r 62000_26000_M1 62000_26000_M2 0.050
r 62000_28000_M1 62000_28000_M2 0.050
r 62000_30000_M1 62000_30000_M2 0.050
r 62000_32000_M1 62000_32000_M2 0.050
r 62000_34000_M1 62000_34000_M2 0.050
r 62000_36000_M1 62000_36000_M2 0.050
r 62000_38000_M1 62000_38000_M2 0.050
r 62000_40000_M1 62000_40000_M2 0.050
r 62000_42000_M1 62000_42000_M2 0.050
r 62000_44000_M1 62000_44000_M2 0.050
r 62000_46000_M1 62000_46000_M2 0.050
r 62000_48000_M1 62000_48000_M2 0.050
r 62000_50000_M1 62000_50000_M2 0.050
r 62000_52000_M1 62000_52000_M2 0.050
r 62000_54000_M1 62000_54000_M2 0.050
r 62000_56000_M1 62000_56000_M2 0.050
r 62000_58000_M1 62000_58000_M2 0.050
r 62000_60000_M1 62000_60000_M2 0.050
r 62000_62000_M1 62000_62000_M2 0.050
r 62000_64000_M1 62000_64000_M2 0.050
r 62000_66000_M1 62000_66000_M2 0.050
r 62000_68000_M1 62000_68000_M2 0.050
r 62000_70000_M1 62000_70000_M2 0.050
r 62000_72000_M1 62000_72000_M2 0.050
r 62000_74000_M1 62000_74000_M2 0.050
r 62000_76000_M1 62000_76000_M2 0.050
r 62000_78000_M1 62000_78000_M2 0.050
r 62000_80000_M1 62000_80000_M2 0.050
r 62000_82000_M1 62000_82000_M2 0.050
r 62000_84000_M1 62000_84000_M2 0.050
r 62000_86000_M1 62000_86000_M2 0.050
r 62000_88000_M1 62000_88000_M2 0.050
r 62000_90000_M1 62000_90000_M2 0.050
r 62000_92000_M1 62000_92000_M2 0.050
r 62000_94000_M1 62000_94000_M2 0.050
r 62000_96000_M1 62000_96000_M2 0.050
r 62000_98000_M1 62000_98000_M2 0.050
r 62000_100000_M1 62000_100000_M2 0.050
r 64000_2000_M1 64000_2000_M2 0.050
r 64000_4000_M1 64000_4000_M2 0.050
r 64000_6000_M1 64000_6000_M2 0.050
r 64000_8000_M1 64000_8000_M2 0.050
r 64000_10000_M1 64000_10000_M2 0.050
r 64000_12000_M1 64000_12000_M2 0.050
r 64000_14000_M1 64000_14000_M2 0.050
r 64000_16000_M1 64000_16000_M2 0.050
r 64000_18000_M1 64000_18000_M2 0.050
r 64000_20000_M1 64000_20000_M2 0.050
r 64000_22000_M1 64000_22000_M2 0.050
r 64000_24000_M1 64000_24000_M2 0.050
r 64000_26000_M1 64000_26000_M2 0.050
r 64000_28000_M1 64000_28000_M2 0.050
r 64000_30000_M1 64000_30000_M2 0.050
r 64000_32000_M1 64000_32000_M2 0.050
r 64000_34000_M1 64000_34000_M2 0.050
r 64000_36000_M1 64000_36000_M2 0.050
r 64000_38000_M1 64000_38000_M2 0.050
r 64000_40000_M1 64000_40000_M2 0.050
r 64000_42000_M1 64000_42000_M2 0.050
r 64000_44000_M1 64000_44000_M2 0.050
r 64000_46000_M1 64000_46000_M2 0.050
r 64000_48000_M1 64000_48000_M2 0.050
r 64000_50000_M1 64000_50000_M2 0.050
r 64000_52000_M1 64000_52000_M2 0.050
r 64000_54000_M1 64000_54000_M2 0.050
r 64000_56000_M1 64000_56000_M2 0.050
r 64000_58000_M1 64000_58000_M2 0.050
r 64000_60000_M1 64000_60000_M2 0.050
r 64000_62000_M1 64000_62000_M2 0.050
r 64000_64000_M1 64000_64000_M2 0.050
r 64000_66000_M1 64000_66000_M2 0.050
r 64000_68000_M1 64000_68000_M2 0.050
r 64000_70000_M1 64000_70000_M2 0.050
r 64000_72000_M1 64000_72000_M2 0.050
r 64000_74000_M1 64000_74000_M2 0.050
r 64000_76000_M1 64000_76000_M2 0.050
r 64000_78000_M1 64000_78000_M2 0.050
r 64000_80000_M1 64000_80000_M2 0.050
r 64000_82000_M1 64000_82000_M2 0.050
r 64000_84000_M1 64000_84000_M2 0.050
r 64000_86000_M1 64000_86000_M2 0.050
r 64000_88000_M1 64000_88000_M2 0.050
r 64000_90000_M1 64000_90000_M2 0.050
r 64000_92000_M1 64000_92000_M2 0.050
r 64000_94000_M1 64000_94000_M2 0.050
r 64000_96000_M1 64000_96000_M2 0.050
r 64000_98000_M1 64000_98000_M2 0.050
r 64000_100000_M1 64000_100000_M2 0.050
r 66000_2000_M1 66000_2000_M2 0.050
r 66000_4000_M1 66000_4000_M2 0.050
r 66000_6000_M1 66000_6000_M2 0.050
r 66000_8000_M1 66000_8000_M2 0.050
r 66000_10000_M1 66000_10000_M2 0.050
r 66000_12000_M1 66000_12000_M2 0.050
r 66000_14000_M1 66000_14000_M2 0.050
r 66000_16000_M1 66000_16000_M2 0.050
r 66000_18000_M1 66000_18000_M2 0.050
r 66000_20000_M1 66000_20000_M2 0.050
r 66000_22000_M1 66000_22000_M2 0.050
r 66000_24000_M1 66000_24000_M2 0.050
r 66000_26000_M1 66000_26000_M2 0.050
r 66000_28000_M1 66000_28000_M2 0.050
r 66000_30000_M1 66000_30000_M2 0.050
r 66000_32000_M1 66000_32000_M2 0.050
r 66000_34000_M1 66000_34000_M2 0.050
r 66000_36000_M1 66000_36000_M2 0.050
r 66000_38000_M1 66000_38000_M2 0.050
r 66000_40000_M1 66000_40000_M2 0.050
r 66000_42000_M1 66000_42000_M2 0.050
r 66000_44000_M1 66000_44000_M2 0.050
r 66000_46000_M1 66000_46000_M2 0.050
r 66000_48000_M1 66000_48000_M2 0.050
r 66000_50000_M1 66000_50000_M2 0.050
r 66000_52000_M1 66000_52000_M2 0.050
r 66000_54000_M1 66000_54000_M2 0.050
r 66000_56000_M1 66000_56000_M2 0.050
r 66000_58000_M1 66000_58000_M2 0.050
r 66000_60000_M1 66000_60000_M2 0.050
r 66000_62000_M1 66000_62000_M2 0.050
r 66000_64000_M1 66000_64000_M2 0.050
r 66000_66000_M1 66000_66000_M2 0.050
r 66000_68000_M1 66000_68000_M2 0.050
r 66000_70000_M1 66000_70000_M2 0.050
r 66000_72000_M1 66000_72000_M2 0.050
r 66000_74000_M1 66000_74000_M2 0.050
r 66000_76000_M1 66000_76000_M2 0.050
r 66000_78000_M1 66000_78000_M2 0.050
r 66000_80000_M1 66000_80000_M2 0.050
r 66000_82000_M1 66000_82000_M2 0.050
r 66000_84000_M1 66000_84000_M2 0.050
r 66000_86000_M1 66000_86000_M2 0.050
r 66000_88000_M1 66000_88000_M2 0.050
r 66000_90000_M1 66000_90000_M2 0.050
r 66000_92000_M1 66000_92000_M2 0.050
r 66000_94000_M1 66000_94000_M2 0.050
r 66000_96000_M1 66000_96000_M2 0.050
r 66000_98000_M1 66000_98000_M2 0.050
r 66000_100000_M1 66000_100000_M2 0.050
r 68000_2000_M1 68000_2000_M2 0.050
r 68000_4000_M1 68000_4000_M2 0.050
r 68000_6000_M1 68000_6000_M2 0.050
r 68000_8000_M1 68000_8000_M2 0.050
r 68000_10000_M1 68000_10000_M2 0.050
r 68000_12000_M1 68000_12000_M2 0.050
r 68000_14000_M1 68000_14000_M2 0.050
r 68000_16000_M1 68000_16000_M2 0.050
r 68000_18000_M1 68000_18000_M2 0.050
r 68000_20000_M1 68000_20000_M2 0.050
r 68000_22000_M1 68000_22000_M2 0.050
r 68000_24000_M1 68000_24000_M2 0.050
r 68000_26000_M1 68000_26000_M2 0.050
r 68000_28000_M1 68000_28000_M2 0.050
r 68000_30000_M1 68000_30000_M2 0.050
r 68000_32000_M1 68000_32000_M2 0.050
r 68000_34000_M1 68000_34000_M2 0.050
r 68000_36000_M1 68000_36000_M2 0.050
r 68000_38000_M1 68000_38000_M2 0.050
r 68000_40000_M1 68000_40000_M2 0.050
r 68000_42000_M1 68000_42000_M2 0.050
r 68000_44000_M1 68000_44000_M2 0.050
r 68000_46000_M1 68000_46000_M2 0.050
r 68000_48000_M1 68000_48000_M2 0.050
r 68000_50000_M1 68000_50000_M2 0.050
r 68000_52000_M1 68000_52000_M2 0.050
r 68000_54000_M1 68000_54000_M2 0.050
r 68000_56000_M1 68000_56000_M2 0.050
r 68000_58000_M1 68000_58000_M2 0.050
r 68000_60000_M1 68000_60000_M2 0.050
r 68000_62000_M1 68000_62000_M2 0.050
r 68000_64000_M1 68000_64000_M2 0.050
r 68000_66000_M1 68000_66000_M2 0.050
r 68000_68000_M1 68000_68000_M2 0.050
r 68000_70000_M1 68000_70000_M2 0.050
r 68000_72000_M1 68000_72000_M2 0.050
r 68000_74000_M1 68000_74000_M2 0.050
r 68000_76000_M1 68000_76000_M2 0.050
r 68000_78000_M1 68000_78000_M2 0.050
r 68000_80000_M1 68000_80000_M2 0.050
r 68000_82000_M1 68000_82000_M2 0.050
r 68000_84000_M1 68000_84000_M2 0.050
r 68000_86000_M1 68000_86000_M2 0.050
r 68000_88000_M1 68000_88000_M2 0.050
r 68000_90000_M1 68000_90000_M2 0.050
r 68000_92000_M1 68000_92000_M2 0.050
r 68000_94000_M1 68000_94000_M2 0.050
r 68000_96000_M1 68000_96000_M2 0.050
r 68000_98000_M1 68000_98000_M2 0.050
r 68000_100000_M1 68000_100000_M2 0.050
r 70000_2000_M1 70000_2000_M2 0.050
r 70000_4000_M1 70000_4000_M2 0.050
r 70000_6000_M1 70000_6000_M2 0.050
r 70000_8000_M1 70000_8000_M2 0.050
r 70000_10000_M1 70000_10000_M2 0.050
r 70000_12000_M1 70000_12000_M2 0.050
r 70000_14000_M1 70000_14000_M2 0.050
r 70000_16000_M1 70000_16000_M2 0.050
r 70000_18000_M1 70000_18000_M2 0.050
r 70000_20000_M1 70000_20000_M2 0.050
r 70000_22000_M1 70000_22000_M2 0.050
r 70000_24000_M1 70000_24000_M2 0.050
r 70000_26000_M1 70000_26000_M2 0.050
r 70000_28000_M1 70000_28000_M2 0.050
r 70000_30000_M1 70000_30000_M2 0.050
r 70000_32000_M1 70000_32000_M2 0.050
r 70000_34000_M1 70000_34000_M2 0.050
r 70000_36000_M1 70000_36000_M2 0.050
r 70000_38000_M1 70000_38000_M2 0.050
r 70000_40000_M1 70000_40000_M2 0.050
r 70000_42000_M1 70000_42000_M2 0.050
r 70000_44000_M1 70000_44000_M2 0.050
r 70000_46000_M1 70000_46000_M2 0.050
r 70000_48000_M1 70000_48000_M2 0.050
r 70000_50000_M1 70000_50000_M2 0.050
r 70000_52000_M1 70000_52000_M2 0.050
r 70000_54000_M1 70000_54000_M2 0.050
r 70000_56000_M1 70000_56000_M2 0.050
r 70000_58000_M1 70000_58000_M2 0.050
r 70000_60000_M1 70000_60000_M2 0.050
r 70000_62000_M1 70000_62000_M2 0.050
r 70000_64000_M1 70000_64000_M2 0.050
r 70000_66000_M1 70000_66000_M2 0.050
r 70000_68000_M1 70000_68000_M2 0.050
r 70000_70000_M1 70000_70000_M2 0.050
r 70000_72000_M1 70000_72000_M2 0.050
r 70000_74000_M1 70000_74000_M2 0.050
r 70000_76000_M1 70000_76000_M2 0.050
r 70000_78000_M1 70000_78000_M2 0.050
r 70000_80000_M1 70000_80000_M2 0.050
r 70000_82000_M1 70000_82000_M2 0.050
r 70000_84000_M1 70000_84000_M2 0.050
r 70000_86000_M1 70000_86000_M2 0.050
r 70000_88000_M1 70000_88000_M2 0.050
r 70000_90000_M1 70000_90000_M2 0.050
r 70000_92000_M1 70000_92000_M2 0.050
r 70000_94000_M1 70000_94000_M2 0.050
r 70000_96000_M1 70000_96000_M2 0.050
r 70000_98000_M1 70000_98000_M2 0.050
r 70000_100000_M1 70000_100000_M2 0.050
r 72000_2000_M1 72000_2000_M2 0.050
r 72000_4000_M1 72000_4000_M2 0.050
r 72000_6000_M1 72000_6000_M2 0.050
r 72000_8000_M1 72000_8000_M2 0.050
r 72000_10000_M1 72000_10000_M2 0.050
r 72000_12000_M1 72000_12000_M2 0.050
r 72000_14000_M1 72000_14000_M2 0.050
r 72000_16000_M1 72000_16000_M2 0.050
r 72000_18000_M1 72000_18000_M2 0.050
r 72000_20000_M1 72000_20000_M2 0.050
r 72000_22000_M1 72000_22000_M2 0.050
r 72000_24000_M1 72000_24000_M2 0.050
r 72000_26000_M1 72000_26000_M2 0.050
r 72000_28000_M1 72000_28000_M2 0.050
r 72000_30000_M1 72000_30000_M2 0.050
r 72000_32000_M1 72000_32000_M2 0.050
r 72000_34000_M1 72000_34000_M2 0.050
r 72000_36000_M1 72000_36000_M2 0.050
r 72000_38000_M1 72000_38000_M2 0.050
r 72000_40000_M1 72000_40000_M2 0.050
r 72000_42000_M1 72000_42000_M2 0.050
r 72000_44000_M1 72000_44000_M2 0.050
r 72000_46000_M1 72000_46000_M2 0.050
r 72000_48000_M1 72000_48000_M2 0.050
r 72000_50000_M1 72000_50000_M2 0.050
r 72000_52000_M1 72000_52000_M2 0.050
r 72000_54000_M1 72000_54000_M2 0.050
r 72000_56000_M1 72000_56000_M2 0.050
r 72000_58000_M1 72000_58000_M2 0.050
r 72000_60000_M1 72000_60000_M2 0.050
r 72000_62000_M1 72000_62000_M2 0.050
r 72000_64000_M1 72000_64000_M2 0.050
r 72000_66000_M1 72000_66000_M2 0.050
r 72000_68000_M1 72000_68000_M2 0.050
r 72000_70000_M1 72000_70000_M2 0.050
r 72000_72000_M1 72000_72000_M2 0.050
r 72000_74000_M1 72000_74000_M2 0.050
r 72000_76000_M1 72000_76000_M2 0.050
r 72000_78000_M1 72000_78000_M2 0.050
r 72000_80000_M1 72000_80000_M2 0.050
r 72000_82000_M1 72000_82000_M2 0.050
r 72000_84000_M1 72000_84000_M2 0.050
r 72000_86000_M1 72000_86000_M2 0.050
r 72000_88000_M1 72000_88000_M2 0.050
r 72000_90000_M1 72000_90000_M2 0.050
r 72000_92000_M1 72000_92000_M2 0.050
r 72000_94000_M1 72000_94000_M2 0.050
r 72000_96000_M1 72000_96000_M2 0.050
r 72000_98000_M1 72000_98000_M2 0.050
r 72000_100000_M1 72000_100000_M2 0.050
r 74000_2000_M1 74000_2000_M2 0.050
r 74000_4000_M1 74000_4000_M2 0.050
r 74000_6000_M1 74000_6000_M2 0.050
r 74000_8000_M1 74000_8000_M2 0.050
r 74000_10000_M1 74000_10000_M2 0.050
r 74000_12000_M1 74000_12000_M2 0.050
r 74000_14000_M1 74000_14000_M2 0.050
r 74000_16000_M1 74000_16000_M2 0.050
r 74000_18000_M1 74000_18000_M2 0.050
r 74000_20000_M1 74000_20000_M2 0.050
r 74000_22000_M1 74000_22000_M2 0.050
r 74000_24000_M1 74000_24000_M2 0.050
r 74000_26000_M1 74000_26000_M2 0.050
r 74000_28000_M1 74000_28000_M2 0.050
r 74000_30000_M1 74000_30000_M2 0.050
r 74000_32000_M1 74000_32000_M2 0.050
r 74000_34000_M1 74000_34000_M2 0.050
r 74000_36000_M1 74000_36000_M2 0.050
r 74000_38000_M1 74000_38000_M2 0.050
r 74000_40000_M1 74000_40000_M2 0.050
r 74000_42000_M1 74000_42000_M2 0.050
r 74000_44000_M1 74000_44000_M2 0.050
r 74000_46000_M1 74000_46000_M2 0.050
r 74000_48000_M1 74000_48000_M2 0.050
r 74000_50000_M1 74000_50000_M2 0.050
r 74000_52000_M1 74000_52000_M2 0.050
r 74000_54000_M1 74000_54000_M2 0.050
r 74000_56000_M1 74000_56000_M2 0.050
r 74000_58000_M1 74000_58000_M2 0.050
r 74000_60000_M1 74000_60000_M2 0.050
r 74000_62000_M1 74000_62000_M2 0.050
r 74000_64000_M1 74000_64000_M2 0.050
r 74000_66000_M1 74000_66000_M2 0.050
r 74000_68000_M1 74000_68000_M2 0.050
r 74000_70000_M1 74000_70000_M2 0.050
r 74000_72000_M1 74000_72000_M2 0.050
r 74000_74000_M1 74000_74000_M2 0.050
r 74000_76000_M1 74000_76000_M2 0.050
r 74000_78000_M1 74000_78000_M2 0.050
r 74000_80000_M1 74000_80000_M2 0.050
r 74000_82000_M1 74000_82000_M2 0.050
r 74000_84000_M1 74000_84000_M2 0.050
r 74000_86000_M1 74000_86000_M2 0.050
r 74000_88000_M1 74000_88000_M2 0.050
r 74000_90000_M1 74000_90000_M2 0.050
r 74000_92000_M1 74000_92000_M2 0.050
r 74000_94000_M1 74000_94000_M2 0.050
r 74000_96000_M1 74000_96000_M2 0.050
r 74000_98000_M1 74000_98000_M2 0.050
r 74000_100000_M1 74000_100000_M2 0.050
r 76000_2000_M1 76000_2000_M2 0.050
r 76000_4000_M1 76000_4000_M2 0.050
r 76000_6000_M1 76000_6000_M2 0.050
r 76000_8000_M1 76000_8000_M2 0.050
r 76000_10000_M1 76000_10000_M2 0.050
r 76000_12000_M1 76000_12000_M2 0.050
r 76000_14000_M1 76000_14000_M2 0.050
r 76000_16000_M1 76000_16000_M2 0.050
r 76000_18000_M1 76000_18000_M2 0.050
r 76000_20000_M1 76000_20000_M2 0.050
r 76000_22000_M1 76000_22000_M2 0.050
r 76000_24000_M1 76000_24000_M2 0.050
r 76000_26000_M1 76000_26000_M2 0.050
r 76000_28000_M1 76000_28000_M2 0.050
r 76000_30000_M1 76000_30000_M2 0.050
r 76000_32000_M1 76000_32000_M2 0.050
r 76000_34000_M1 76000_34000_M2 0.050
r 76000_36000_M1 76000_36000_M2 0.050
r 76000_38000_M1 76000_38000_M2 0.050
r 76000_40000_M1 76000_40000_M2 0.050
r 76000_42000_M1 76000_42000_M2 0.050
r 76000_44000_M1 76000_44000_M2 0.050
r 76000_46000_M1 76000_46000_M2 0.050
r 76000_48000_M1 76000_48000_M2 0.050
r 76000_50000_M1 76000_50000_M2 0.050
r 76000_52000_M1 76000_52000_M2 0.050
r 76000_54000_M1 76000_54000_M2 0.050
r 76000_56000_M1 76000_56000_M2 0.050
r 76000_58000_M1 76000_58000_M2 0.050
r 76000_60000_M1 76000_60000_M2 0.050
r 76000_62000_M1 76000_62000_M2 0.050
r 76000_64000_M1 76000_64000_M2 0.050
r 76000_66000_M1 76000_66000_M2 0.050
r 76000_68000_M1 76000_68000_M2 0.050
r 76000_70000_M1 76000_70000_M2 0.050
r 76000_72000_M1 76000_72000_M2 0.050
r 76000_74000_M1 76000_74000_M2 0.050
r 76000_76000_M1 76000_76000_M2 0.050
r 76000_78000_M1 76000_78000_M2 0.050
r 76000_80000_M1 76000_80000_M2 0.050
r 76000_82000_M1 76000_82000_M2 0.050
r 76000_84000_M1 76000_84000_M2 0.050
r 76000_86000_M1 76000_86000_M2 0.050
r 76000_88000_M1 76000_88000_M2 0.050
r 76000_90000_M1 76000_90000_M2 0.050
r 76000_92000_M1 76000_92000_M2 0.050
r 76000_94000_M1 76000_94000_M2 0.050
r 76000_96000_M1 76000_96000_M2 0.050
r 76000_98000_M1 76000_98000_M2 0.050
r 76000_100000_M1 76000_100000_M2 0.050
r 78000_2000_M1 78000_2000_M2 0.050
r 78000_4000_M1 78000_4000_M2 0.050
r 78000_6000_M1 78000_6000_M2 0.050
r 78000_8000_M1 78000_8000_M2 0.050
r 78000_10000_M1 78000_10000_M2 0.050
r 78000_12000_M1 78000_12000_M2 0.050
r 78000_14000_M1 78000_14000_M2 0.050
r 78000_16000_M1 78000_16000_M2 0.050
r 78000_18000_M1 78000_18000_M2 0.050
r 78000_20000_M1 78000_20000_M2 0.050
r 78000_22000_M1 78000_22000_M2 0.050
r 78000_24000_M1 78000_24000_M2 0.050
r 78000_26000_M1 78000_26000_M2 0.050
r 78000_28000_M1 78000_28000_M2 0.050
r 78000_30000_M1 78000_30000_M2 0.050
r 78000_32000_M1 78000_32000_M2 0.050
r 78000_34000_M1 78000_34000_M2 0.050
r 78000_36000_M1 78000_36000_M2 0.050
r 78000_38000_M1 78000_38000_M2 0.050
r 78000_40000_M1 78000_40000_M2 0.050
r 78000_42000_M1 78000_42000_M2 0.050
r 78000_44000_M1 78000_44000_M2 0.050
r 78000_46000_M1 78000_46000_M2 0.050
r 78000_48000_M1 78000_48000_M2 0.050
r 78000_50000_M1 78000_50000_M2 0.050
r 78000_52000_M1 78000_52000_M2 0.050
r 78000_54000_M1 78000_54000_M2 0.050
r 78000_56000_M1 78000_56000_M2 0.050
r 78000_58000_M1 78000_58000_M2 0.050
r 78000_60000_M1 78000_60000_M2 0.050
r 78000_62000_M1 78000_62000_M2 0.050
r 78000_64000_M1 78000_64000_M2 0.050
r 78000_66000_M1 78000_66000_M2 0.050
r 78000_68000_M1 78000_68000_M2 0.050
r 78000_70000_M1 78000_70000_M2 0.050
r 78000_72000_M1 78000_72000_M2 0.050
r 78000_74000_M1 78000_74000_M2 0.050
r 78000_76000_M1 78000_76000_M2 0.050
r 78000_78000_M1 78000_78000_M2 0.050
r 78000_80000_M1 78000_80000_M2 0.050
r 78000_82000_M1 78000_82000_M2 0.050
r 78000_84000_M1 78000_84000_M2 0.050
r 78000_86000_M1 78000_86000_M2 0.050
r 78000_88000_M1 78000_88000_M2 0.050
r 78000_90000_M1 78000_90000_M2 0.050
r 78000_92000_M1 78000_92000_M2 0.050
r 78000_94000_M1 78000_94000_M2 0.050
r 78000_96000_M1 78000_96000_M2 0.050
r 78000_98000_M1 78000_98000_M2 0.050
r 78000_100000_M1 78000_100000_M2 0.050
r 80000_2000_M1 80000_2000_M2 0.050
r 80000_4000_M1 80000_4000_M2 0.050
r 80000_6000_M1 80000_6000_M2 0.050
r 80000_8000_M1 80000_8000_M2 0.050
r 80000_10000_M1 80000_10000_M2 0.050
r 80000_12000_M1 80000_12000_M2 0.050
r 80000_14000_M1 80000_14000_M2 0.050
r 80000_16000_M1 80000_16000_M2 0.050
r 80000_18000_M1 80000_18000_M2 0.050
r 80000_20000_M1 80000_20000_M2 0.050
r 80000_22000_M1 80000_22000_M2 0.050
r 80000_24000_M1 80000_24000_M2 0.050
r 80000_26000_M1 80000_26000_M2 0.050
r 80000_28000_M1 80000_28000_M2 0.050
r 80000_30000_M1 80000_30000_M2 0.050
r 80000_32000_M1 80000_32000_M2 0.050
r 80000_34000_M1 80000_34000_M2 0.050
r 80000_36000_M1 80000_36000_M2 0.050
r 80000_38000_M1 80000_38000_M2 0.050
r 80000_40000_M1 80000_40000_M2 0.050
r 80000_42000_M1 80000_42000_M2 0.050
r 80000_44000_M1 80000_44000_M2 0.050
r 80000_46000_M1 80000_46000_M2 0.050
r 80000_48000_M1 80000_48000_M2 0.050
r 80000_50000_M1 80000_50000_M2 0.050
r 80000_52000_M1 80000_52000_M2 0.050
r 80000_54000_M1 80000_54000_M2 0.050
r 80000_56000_M1 80000_56000_M2 0.050
r 80000_58000_M1 80000_58000_M2 0.050
r 80000_60000_M1 80000_60000_M2 0.050
r 80000_62000_M1 80000_62000_M2 0.050
r 80000_64000_M1 80000_64000_M2 0.050
r 80000_66000_M1 80000_66000_M2 0.050
r 80000_68000_M1 80000_68000_M2 0.050
r 80000_70000_M1 80000_70000_M2 0.050
r 80000_72000_M1 80000_72000_M2 0.050
r 80000_74000_M1 80000_74000_M2 0.050
r 80000_76000_M1 80000_76000_M2 0.050
r 80000_78000_M1 80000_78000_M2 0.050
r 80000_80000_M1 80000_80000_M2 0.050
r 80000_82000_M1 80000_82000_M2 0.050
r 80000_84000_M1 80000_84000_M2 0.050
r 80000_86000_M1 80000_86000_M2 0.050
r 80000_88000_M1 80000_88000_M2 0.050
r 80000_90000_M1 80000_90000_M2 0.050
r 80000_92000_M1 80000_92000_M2 0.050
r 80000_94000_M1 80000_94000_M2 0.050
r 80000_96000_M1 80000_96000_M2 0.050
r 80000_98000_M1 80000_98000_M2 0.050
r 80000_100000_M1 80000_100000_M2 0.050
r 82000_2000_M1 82000_2000_M2 0.050
r 82000_4000_M1 82000_4000_M2 0.050
r 82000_6000_M1 82000_6000_M2 0.050
r 82000_8000_M1 82000_8000_M2 0.050
r 82000_10000_M1 82000_10000_M2 0.050
r 82000_12000_M1 82000_12000_M2 0.050
r 82000_14000_M1 82000_14000_M2 0.050
r 82000_16000_M1 82000_16000_M2 0.050
r 82000_18000_M1 82000_18000_M2 0.050
r 82000_20000_M1 82000_20000_M2 0.050
r 82000_22000_M1 82000_22000_M2 0.050
r 82000_24000_M1 82000_24000_M2 0.050
r 82000_26000_M1 82000_26000_M2 0.050
r 82000_28000_M1 82000_28000_M2 0.050
r 82000_30000_M1 82000_30000_M2 0.050
r 82000_32000_M1 82000_32000_M2 0.050
r 82000_34000_M1 82000_34000_M2 0.050
r 82000_36000_M1 82000_36000_M2 0.050
r 82000_38000_M1 82000_38000_M2 0.050
r 82000_40000_M1 82000_40000_M2 0.050
r 82000_42000_M1 82000_42000_M2 0.050
r 82000_44000_M1 82000_44000_M2 0.050
r 82000_46000_M1 82000_46000_M2 0.050
r 82000_48000_M1 82000_48000_M2 0.050
r 82000_50000_M1 82000_50000_M2 0.050
r 82000_52000_M1 82000_52000_M2 0.050
r 82000_54000_M1 82000_54000_M2 0.050
r 82000_56000_M1 82000_56000_M2 0.050
r 82000_58000_M1 82000_58000_M2 0.050
r 82000_60000_M1 82000_60000_M2 0.050
r 82000_62000_M1 82000_62000_M2 0.050
r 82000_64000_M1 82000_64000_M2 0.050
r 82000_66000_M1 82000_66000_M2 0.050
r 82000_68000_M1 82000_68000_M2 0.050
r 82000_70000_M1 82000_70000_M2 0.050
r 82000_72000_M1 82000_72000_M2 0.050
r 82000_74000_M1 82000_74000_M2 0.050
r 82000_76000_M1 82000_76000_M2 0.050
r 82000_78000_M1 82000_78000_M2 0.050
r 82000_80000_M1 82000_80000_M2 0.050
r 82000_82000_M1 82000_82000_M2 0.050
r 82000_84000_M1 82000_84000_M2 0.050
r 82000_86000_M1 82000_86000_M2 0.050
r 82000_88000_M1 82000_88000_M2 0.050
r 82000_90000_M1 82000_90000_M2 0.050
r 82000_92000_M1 82000_92000_M2 0.050
r 82000_94000_M1 82000_94000_M2 0.050
r 82000_96000_M1 82000_96000_M2 0.050
r 82000_98000_M1 82000_98000_M2 0.050
r 82000_100000_M1 82000_100000_M2 0.050
r 84000_2000_M1 84000_2000_M2 0.050
r 84000_4000_M1 84000_4000_M2 0.050
r 84000_6000_M1 84000_6000_M2 0.050
r 84000_8000_M1 84000_8000_M2 0.050
r 84000_10000_M1 84000_10000_M2 0.050
r 84000_12000_M1 84000_12000_M2 0.050
r 84000_14000_M1 84000_14000_M2 0.050
r 84000_16000_M1 84000_16000_M2 0.050
r 84000_18000_M1 84000_18000_M2 0.050
r 84000_20000_M1 84000_20000_M2 0.050
r 84000_22000_M1 84000_22000_M2 0.050
r 84000_24000_M1 84000_24000_M2 0.050
r 84000_26000_M1 84000_26000_M2 0.050
r 84000_28000_M1 84000_28000_M2 0.050
r 84000_30000_M1 84000_30000_M2 0.050
r 84000_32000_M1 84000_32000_M2 0.050
r 84000_34000_M1 84000_34000_M2 0.050
r 84000_36000_M1 84000_36000_M2 0.050
r 84000_38000_M1 84000_38000_M2 0.050
r 84000_40000_M1 84000_40000_M2 0.050
r 84000_42000_M1 84000_42000_M2 0.050
r 84000_44000_M1 84000_44000_M2 0.050
r 84000_46000_M1 84000_46000_M2 0.050
r 84000_48000_M1 84000_48000_M2 0.050
r 84000_50000_M1 84000_50000_M2 0.050
r 84000_52000_M1 84000_52000_M2 0.050
r 84000_54000_M1 84000_54000_M2 0.050
r 84000_56000_M1 84000_56000_M2 0.050
r 84000_58000_M1 84000_58000_M2 0.050
r 84000_60000_M1 84000_60000_M2 0.050
r 84000_62000_M1 84000_62000_M2 0.050
r 84000_64000_M1 84000_64000_M2 0.050
r 84000_66000_M1 84000_66000_M2 0.050
r 84000_68000_M1 84000_68000_M2 0.050
r 84000_70000_M1 84000_70000_M2 0.050
r 84000_72000_M1 84000_72000_M2 0.050
r 84000_74000_M1 84000_74000_M2 0.050
r 84000_76000_M1 84000_76000_M2 0.050
r 84000_78000_M1 84000_78000_M2 0.050
r 84000_80000_M1 84000_80000_M2 0.050
r 84000_82000_M1 84000_82000_M2 0.050
r 84000_84000_M1 84000_84000_M2 0.050
r 84000_86000_M1 84000_86000_M2 0.050
r 84000_88000_M1 84000_88000_M2 0.050
r 84000_90000_M1 84000_90000_M2 0.050
r 84000_92000_M1 84000_92000_M2 0.050
r 84000_94000_M1 84000_94000_M2 0.050
r 84000_96000_M1 84000_96000_M2 0.050
r 84000_98000_M1 84000_98000_M2 0.050
r 84000_100000_M1 84000_100000_M2 0.050
r 86000_2000_M1 86000_2000_M2 0.050
r 86000_4000_M1 86000_4000_M2 0.050
r 86000_6000_M1 86000_6000_M2 0.050
r 86000_8000_M1 86000_8000_M2 0.050
r 86000_10000_M1 86000_10000_M2 0.050
r 86000_12000_M1 86000_12000_M2 0.050
r 86000_14000_M1 86000_14000_M2 0.050
r 86000_16000_M1 86000_16000_M2 0.050
r 86000_18000_M1 86000_18000_M2 0.050
r 86000_20000_M1 86000_20000_M2 0.050
r 86000_22000_M1 86000_22000_M2 0.050
r 86000_24000_M1 86000_24000_M2 0.050
r 86000_26000_M1 86000_26000_M2 0.050
r 86000_28000_M1 86000_28000_M2 0.050
r 86000_30000_M1 86000_30000_M2 0.050
r 86000_32000_M1 86000_32000_M2 0.050
r 86000_34000_M1 86000_34000_M2 0.050
r 86000_36000_M1 86000_36000_M2 0.050
r 86000_38000_M1 86000_38000_M2 0.050
r 86000_40000_M1 86000_40000_M2 0.050
r 86000_42000_M1 86000_42000_M2 0.050
r 86000_44000_M1 86000_44000_M2 0.050
r 86000_46000_M1 86000_46000_M2 0.050
r 86000_48000_M1 86000_48000_M2 0.050
r 86000_50000_M1 86000_50000_M2 0.050
r 86000_52000_M1 86000_52000_M2 0.050
r 86000_54000_M1 86000_54000_M2 0.050
r 86000_56000_M1 86000_56000_M2 0.050
r 86000_58000_M1 86000_58000_M2 0.050
r 86000_60000_M1 86000_60000_M2 0.050
r 86000_62000_M1 86000_62000_M2 0.050
r 86000_64000_M1 86000_64000_M2 0.050
r 86000_66000_M1 86000_66000_M2 0.050
r 86000_68000_M1 86000_68000_M2 0.050
r 86000_70000_M1 86000_70000_M2 0.050
r 86000_72000_M1 86000_72000_M2 0.050
r 86000_74000_M1 86000_74000_M2 0.050
r 86000_76000_M1 86000_76000_M2 0.050
r 86000_78000_M1 86000_78000_M2 0.050
r 86000_80000_M1 86000_80000_M2 0.050
r 86000_82000_M1 86000_82000_M2 0.050
r 86000_84000_M1 86000_84000_M2 0.050
r 86000_86000_M1 86000_86000_M2 0.050
r 86000_88000_M1 86000_88000_M2 0.050
r 86000_90000_M1 86000_90000_M2 0.050
r 86000_92000_M1 86000_92000_M2 0.050
r 86000_94000_M1 86000_94000_M2 0.050
r 86000_96000_M1 86000_96000_M2 0.050
r 86000_98000_M1 86000_98000_M2 0.050
r 86000_100000_M1 86000_100000_M2 0.050
r 88000_2000_M1 88000_2000_M2 0.050
r 88000_4000_M1 88000_4000_M2 0.050
r 88000_6000_M1 88000_6000_M2 0.050
r 88000_8000_M1 88000_8000_M2 0.050
r 88000_10000_M1 88000_10000_M2 0.050
r 88000_12000_M1 88000_12000_M2 0.050
r 88000_14000_M1 88000_14000_M2 0.050
r 88000_16000_M1 88000_16000_M2 0.050
r 88000_18000_M1 88000_18000_M2 0.050
r 88000_20000_M1 88000_20000_M2 0.050
r 88000_22000_M1 88000_22000_M2 0.050
r 88000_24000_M1 88000_24000_M2 0.050
r 88000_26000_M1 88000_26000_M2 0.050
r 88000_28000_M1 88000_28000_M2 0.050
r 88000_30000_M1 88000_30000_M2 0.050
r 88000_32000_M1 88000_32000_M2 0.050
r 88000_34000_M1 88000_34000_M2 0.050
r 88000_36000_M1 88000_36000_M2 0.050
r 88000_38000_M1 88000_38000_M2 0.050
r 88000_40000_M1 88000_40000_M2 0.050
r 88000_42000_M1 88000_42000_M2 0.050
r 88000_44000_M1 88000_44000_M2 0.050
r 88000_46000_M1 88000_46000_M2 0.050
r 88000_48000_M1 88000_48000_M2 0.050
r 88000_50000_M1 88000_50000_M2 0.050
r 88000_52000_M1 88000_52000_M2 0.050
r 88000_54000_M1 88000_54000_M2 0.050
r 88000_56000_M1 88000_56000_M2 0.050
r 88000_58000_M1 88000_58000_M2 0.050
r 88000_60000_M1 88000_60000_M2 0.050
r 88000_62000_M1 88000_62000_M2 0.050
r 88000_64000_M1 88000_64000_M2 0.050
r 88000_66000_M1 88000_66000_M2 0.050
r 88000_68000_M1 88000_68000_M2 0.050
r 88000_70000_M1 88000_70000_M2 0.050
r 88000_72000_M1 88000_72000_M2 0.050
r 88000_74000_M1 88000_74000_M2 0.050
r 88000_76000_M1 88000_76000_M2 0.050
r 88000_78000_M1 88000_78000_M2 0.050
r 88000_80000_M1 88000_80000_M2 0.050
r 88000_82000_M1 88000_82000_M2 0.050
r 88000_84000_M1 88000_84000_M2 0.050
r 88000_86000_M1 88000_86000_M2 0.050
r 88000_88000_M1 88000_88000_M2 0.050
r 88000_90000_M1 88000_90000_M2 0.050
r 88000_92000_M1 88000_92000_M2 0.050
r 88000_94000_M1 88000_94000_M2 0.050
r 88000_96000_M1 88000_96000_M2 0.050
r 88000_98000_M1 88000_98000_M2 0.050
r 88000_100000_M1 88000_100000_M2 0.050
r 90000_2000_M1 90000_2000_M2 0.050
r 90000_4000_M1 90000_4000_M2 0.050
r 90000_6000_M1 90000_6000_M2 0.050
r 90000_8000_M1 90000_8000_M2 0.050
r 90000_10000_M1 90000_10000_M2 0.050
r 90000_12000_M1 90000_12000_M2 0.050
r 90000_14000_M1 90000_14000_M2 0.050
r 90000_16000_M1 90000_16000_M2 0.050
r 90000_18000_M1 90000_18000_M2 0.050
r 90000_20000_M1 90000_20000_M2 0.050
r 90000_22000_M1 90000_22000_M2 0.050
r 90000_24000_M1 90000_24000_M2 0.050
r 90000_26000_M1 90000_26000_M2 0.050
r 90000_28000_M1 90000_28000_M2 0.050
r 90000_30000_M1 90000_30000_M2 0.050
r 90000_32000_M1 90000_32000_M2 0.050
r 90000_34000_M1 90000_34000_M2 0.050
r 90000_36000_M1 90000_36000_M2 0.050
r 90000_38000_M1 90000_38000_M2 0.050
r 90000_40000_M1 90000_40000_M2 0.050
r 90000_42000_M1 90000_42000_M2 0.050
r 90000_44000_M1 90000_44000_M2 0.050
r 90000_46000_M1 90000_46000_M2 0.050
r 90000_48000_M1 90000_48000_M2 0.050
r 90000_50000_M1 90000_50000_M2 0.050
r 90000_52000_M1 90000_52000_M2 0.050
r 90000_54000_M1 90000_54000_M2 0.050
r 90000_56000_M1 90000_56000_M2 0.050
r 90000_58000_M1 90000_58000_M2 0.050
r 90000_60000_M1 90000_60000_M2 0.050
r 90000_62000_M1 90000_62000_M2 0.050
r 90000_64000_M1 90000_64000_M2 0.050
r 90000_66000_M1 90000_66000_M2 0.050
r 90000_68000_M1 90000_68000_M2 0.050
r 90000_70000_M1 90000_70000_M2 0.050
r 90000_72000_M1 90000_72000_M2 0.050
r 90000_74000_M1 90000_74000_M2 0.050
r 90000_76000_M1 90000_76000_M2 0.050
r 90000_78000_M1 90000_78000_M2 0.050
r 90000_80000_M1 90000_80000_M2 0.050
r 90000_82000_M1 90000_82000_M2 0.050
r 90000_84000_M1 90000_84000_M2 0.050
r 90000_86000_M1 90000_86000_M2 0.050
r 90000_88000_M1 90000_88000_M2 0.050
r 90000_90000_M1 90000_90000_M2 0.050
r 90000_92000_M1 90000_92000_M2 0.050
r 90000_94000_M1 90000_94000_M2 0.050
r 90000_96000_M1 90000_96000_M2 0.050
r 90000_98000_M1 90000_98000_M2 0.050
r 90000_100000_M1 90000_100000_M2 0.050
r 92000_2000_M1 92000_2000_M2 0.050
r 92000_4000_M1 92000_4000_M2 0.050
r 92000_6000_M1 92000_6000_M2 0.050
r 92000_8000_M1 92000_8000_M2 0.050
r 92000_10000_M1 92000_10000_M2 0.050
r 92000_12000_M1 92000_12000_M2 0.050
r 92000_14000_M1 92000_14000_M2 0.050
r 92000_16000_M1 92000_16000_M2 0.050
r 92000_18000_M1 92000_18000_M2 0.050
r 92000_20000_M1 92000_20000_M2 0.050
r 92000_22000_M1 92000_22000_M2 0.050
r 92000_24000_M1 92000_24000_M2 0.050
r 92000_26000_M1 92000_26000_M2 0.050
r 92000_28000_M1 92000_28000_M2 0.050
r 92000_30000_M1 92000_30000_M2 0.050
r 92000_32000_M1 92000_32000_M2 0.050
r 92000_34000_M1 92000_34000_M2 0.050
r 92000_36000_M1 92000_36000_M2 0.050
r 92000_38000_M1 92000_38000_M2 0.050
r 92000_40000_M1 92000_40000_M2 0.050
r 92000_42000_M1 92000_42000_M2 0.050
r 92000_44000_M1 92000_44000_M2 0.050
r 92000_46000_M1 92000_46000_M2 0.050
r 92000_48000_M1 92000_48000_M2 0.050
r 92000_50000_M1 92000_50000_M2 0.050
r 92000_52000_M1 92000_52000_M2 0.050
r 92000_54000_M1 92000_54000_M2 0.050
r 92000_56000_M1 92000_56000_M2 0.050
r 92000_58000_M1 92000_58000_M2 0.050
r 92000_60000_M1 92000_60000_M2 0.050
r 92000_62000_M1 92000_62000_M2 0.050
r 92000_64000_M1 92000_64000_M2 0.050
r 92000_66000_M1 92000_66000_M2 0.050
r 92000_68000_M1 92000_68000_M2 0.050
r 92000_70000_M1 92000_70000_M2 0.050
r 92000_72000_M1 92000_72000_M2 0.050
r 92000_74000_M1 92000_74000_M2 0.050
r 92000_76000_M1 92000_76000_M2 0.050
r 92000_78000_M1 92000_78000_M2 0.050
r 92000_80000_M1 92000_80000_M2 0.050
r 92000_82000_M1 92000_82000_M2 0.050
r 92000_84000_M1 92000_84000_M2 0.050
r 92000_86000_M1 92000_86000_M2 0.050
r 92000_88000_M1 92000_88000_M2 0.050
r 92000_90000_M1 92000_90000_M2 0.050
r 92000_92000_M1 92000_92000_M2 0.050
r 92000_94000_M1 92000_94000_M2 0.050
r 92000_96000_M1 92000_96000_M2 0.050
r 92000_98000_M1 92000_98000_M2 0.050
r 92000_100000_M1 92000_100000_M2 0.050
r 94000_2000_M1 94000_2000_M2 0.050
r 94000_4000_M1 94000_4000_M2 0.050
r 94000_6000_M1 94000_6000_M2 0.050
r 94000_8000_M1 94000_8000_M2 0.050
r 94000_10000_M1 94000_10000_M2 0.050
r 94000_12000_M1 94000_12000_M2 0.050
r 94000_14000_M1 94000_14000_M2 0.050
r 94000_16000_M1 94000_16000_M2 0.050
r 94000_18000_M1 94000_18000_M2 0.050
r 94000_20000_M1 94000_20000_M2 0.050
r 94000_22000_M1 94000_22000_M2 0.050
r 94000_24000_M1 94000_24000_M2 0.050
r 94000_26000_M1 94000_26000_M2 0.050
r 94000_28000_M1 94000_28000_M2 0.050
r 94000_30000_M1 94000_30000_M2 0.050
r 94000_32000_M1 94000_32000_M2 0.050
r 94000_34000_M1 94000_34000_M2 0.050
r 94000_36000_M1 94000_36000_M2 0.050
r 94000_38000_M1 94000_38000_M2 0.050
r 94000_40000_M1 94000_40000_M2 0.050
r 94000_42000_M1 94000_42000_M2 0.050
r 94000_44000_M1 94000_44000_M2 0.050
r 94000_46000_M1 94000_46000_M2 0.050
r 94000_48000_M1 94000_48000_M2 0.050
r 94000_50000_M1 94000_50000_M2 0.050
r 94000_52000_M1 94000_52000_M2 0.050
r 94000_54000_M1 94000_54000_M2 0.050
r 94000_56000_M1 94000_56000_M2 0.050
r 94000_58000_M1 94000_58000_M2 0.050
r 94000_60000_M1 94000_60000_M2 0.050
r 94000_62000_M1 94000_62000_M2 0.050
r 94000_64000_M1 94000_64000_M2 0.050
r 94000_66000_M1 94000_66000_M2 0.050
r 94000_68000_M1 94000_68000_M2 0.050
r 94000_70000_M1 94000_70000_M2 0.050
r 94000_72000_M1 94000_72000_M2 0.050
r 94000_74000_M1 94000_74000_M2 0.050
r 94000_76000_M1 94000_76000_M2 0.050
r 94000_78000_M1 94000_78000_M2 0.050
r 94000_80000_M1 94000_80000_M2 0.050
r 94000_82000_M1 94000_82000_M2 0.050
r 94000_84000_M1 94000_84000_M2 0.050
r 94000_86000_M1 94000_86000_M2 0.050
r 94000_88000_M1 94000_88000_M2 0.050
r 94000_90000_M1 94000_90000_M2 0.050
r 94000_92000_M1 94000_92000_M2 0.050
r 94000_94000_M1 94000_94000_M2 0.050
r 94000_96000_M1 94000_96000_M2 0.050
r 94000_98000_M1 94000_98000_M2 0.050
r 94000_100000_M1 94000_100000_M2 0.050
r 96000_2000_M1 96000_2000_M2 0.050
r 96000_4000_M1 96000_4000_M2 0.050
r 96000_6000_M1 96000_6000_M2 0.050
r 96000_8000_M1 96000_8000_M2 0.050
r 96000_10000_M1 96000_10000_M2 0.050
r 96000_12000_M1 96000_12000_M2 0.050
r 96000_14000_M1 96000_14000_M2 0.050
r 96000_16000_M1 96000_16000_M2 0.050
r 96000_18000_M1 96000_18000_M2 0.050
r 96000_20000_M1 96000_20000_M2 0.050
r 96000_22000_M1 96000_22000_M2 0.050
r 96000_24000_M1 96000_24000_M2 0.050
r 96000_26000_M1 96000_26000_M2 0.050
r 96000_28000_M1 96000_28000_M2 0.050
r 96000_30000_M1 96000_30000_M2 0.050
r 96000_32000_M1 96000_32000_M2 0.050
r 96000_34000_M1 96000_34000_M2 0.050
r 96000_36000_M1 96000_36000_M2 0.050
r 96000_38000_M1 96000_38000_M2 0.050
r 96000_40000_M1 96000_40000_M2 0.050
r 96000_42000_M1 96000_42000_M2 0.050
r 96000_44000_M1 96000_44000_M2 0.050
r 96000_46000_M1 96000_46000_M2 0.050
r 96000_48000_M1 96000_48000_M2 0.050
r 96000_50000_M1 96000_50000_M2 0.050
r 96000_52000_M1 96000_52000_M2 0.050
r 96000_54000_M1 96000_54000_M2 0.050
r 96000_56000_M1 96000_56000_M2 0.050
r 96000_58000_M1 96000_58000_M2 0.050
r 96000_60000_M1 96000_60000_M2 0.050
r 96000_62000_M1 96000_62000_M2 0.050
r 96000_64000_M1 96000_64000_M2 0.050
r 96000_66000_M1 96000_66000_M2 0.050
r 96000_68000_M1 96000_68000_M2 0.050
r 96000_70000_M1 96000_70000_M2 0.050
r 96000_72000_M1 96000_72000_M2 0.050
r 96000_74000_M1 96000_74000_M2 0.050
r 96000_76000_M1 96000_76000_M2 0.050
r 96000_78000_M1 96000_78000_M2 0.050
r 96000_80000_M1 96000_80000_M2 0.050
r 96000_82000_M1 96000_82000_M2 0.050
r 96000_84000_M1 96000_84000_M2 0.050
r 96000_86000_M1 96000_86000_M2 0.050
r 96000_88000_M1 96000_88000_M2 0.050
r 96000_90000_M1 96000_90000_M2 0.050
r 96000_92000_M1 96000_92000_M2 0.050
r 96000_94000_M1 96000_94000_M2 0.050
r 96000_96000_M1 96000_96000_M2 0.050
r 96000_98000_M1 96000_98000_M2 0.050
r 96000_100000_M1 96000_100000_M2 0.050
r 98000_2000_M1 98000_2000_M2 0.050
r 98000_4000_M1 98000_4000_M2 0.050
r 98000_6000_M1 98000_6000_M2 0.050
r 98000_8000_M1 98000_8000_M2 0.050
r 98000_10000_M1 98000_10000_M2 0.050
r 98000_12000_M1 98000_12000_M2 0.050
r 98000_14000_M1 98000_14000_M2 0.050
r 98000_16000_M1 98000_16000_M2 0.050
r 98000_18000_M1 98000_18000_M2 0.050
r 98000_20000_M1 98000_20000_M2 0.050
r 98000_22000_M1 98000_22000_M2 0.050
r 98000_24000_M1 98000_24000_M2 0.050
r 98000_26000_M1 98000_26000_M2 0.050
r 98000_28000_M1 98000_28000_M2 0.050
r 98000_30000_M1 98000_30000_M2 0.050
r 98000_32000_M1 98000_32000_M2 0.050
r 98000_34000_M1 98000_34000_M2 0.050
r 98000_36000_M1 98000_36000_M2 0.050
r 98000_38000_M1 98000_38000_M2 0.050
r 98000_40000_M1 98000_40000_M2 0.050
r 98000_42000_M1 98000_42000_M2 0.050
r 98000_44000_M1 98000_44000_M2 0.050
r 98000_46000_M1 98000_46000_M2 0.050
r 98000_48000_M1 98000_48000_M2 0.050
r 98000_50000_M1 98000_50000_M2 0.050
r 98000_52000_M1 98000_52000_M2 0.050
r 98000_54000_M1 98000_54000_M2 0.050
r 98000_56000_M1 98000_56000_M2 0.050
r 98000_58000_M1 98000_58000_M2 0.050
r 98000_60000_M1 98000_60000_M2 0.050
r 98000_62000_M1 98000_62000_M2 0.050
r 98000_64000_M1 98000_64000_M2 0.050
r 98000_66000_M1 98000_66000_M2 0.050
r 98000_68000_M1 98000_68000_M2 0.050
r 98000_70000_M1 98000_70000_M2 0.050
r 98000_72000_M1 98000_72000_M2 0.050
r 98000_74000_M1 98000_74000_M2 0.050
r 98000_76000_M1 98000_76000_M2 0.050
r 98000_78000_M1 98000_78000_M2 0.050
r 98000_80000_M1 98000_80000_M2 0.050
r 98000_82000_M1 98000_82000_M2 0.050
r 98000_84000_M1 98000_84000_M2 0.050
r 98000_86000_M1 98000_86000_M2 0.050
r 98000_88000_M1 98000_88000_M2 0.050
r 98000_90000_M1 98000_90000_M2 0.050
r 98000_92000_M1 98000_92000_M2 0.050
r 98000_94000_M1 98000_94000_M2 0.050
r 98000_96000_M1 98000_96000_M2 0.050
r 98000_98000_M1 98000_98000_M2 0.050
r 98000_100000_M1 98000_100000_M2 0.050
r 100000_2000_M1 100000_2000_M2 0.050
r 100000_4000_M1 100000_4000_M2 0.050
r 100000_6000_M1 100000_6000_M2 0.050
r 100000_8000_M1 100000_8000_M2 0.050
r 100000_10000_M1 100000_10000_M2 0.050
r 100000_12000_M1 100000_12000_M2 0.050
r 100000_14000_M1 100000_14000_M2 0.050
r 100000_16000_M1 100000_16000_M2 0.050
r 100000_18000_M1 100000_18000_M2 0.050
r 100000_20000_M1 100000_20000_M2 0.050
r 100000_22000_M1 100000_22000_M2 0.050
r 100000_24000_M1 100000_24000_M2 0.050
r 100000_26000_M1 100000_26000_M2 0.050
r 100000_28000_M1 100000_28000_M2 0.050
r 100000_30000_M1 100000_30000_M2 0.050
r 100000_32000_M1 100000_32000_M2 0.050
r 100000_34000_M1 100000_34000_M2 0.050
r 100000_36000_M1 100000_36000_M2 0.050
r 100000_38000_M1 100000_38000_M2 0.050
r 100000_40000_M1 100000_40000_M2 0.050
r 100000_42000_M1 100000_42000_M2 0.050
r 100000_44000_M1 100000_44000_M2 0.050
r 100000_46000_M1 100000_46000_M2 0.050
r 100000_48000_M1 100000_48000_M2 0.050
r 100000_50000_M1 100000_50000_M2 0.050
r 100000_52000_M1 100000_52000_M2 0.050
r 100000_54000_M1 100000_54000_M2 0.050
r 100000_56000_M1 100000_56000_M2 0.050
r 100000_58000_M1 100000_58000_M2 0.050
r 100000_60000_M1 100000_60000_M2 0.050
r 100000_62000_M1 100000_62000_M2 0.050
r 100000_64000_M1 100000_64000_M2 0.050
r 100000_66000_M1 100000_66000_M2 0.050
r 100000_68000_M1 100000_68000_M2 0.050
r 100000_70000_M1 100000_70000_M2 0.050
r 100000_72000_M1 100000_72000_M2 0.050
r 100000_74000_M1 100000_74000_M2 0.050
r 100000_76000_M1 100000_76000_M2 0.050
r 100000_78000_M1 100000_78000_M2 0.050
r 100000_80000_M1 100000_80000_M2 0.050
r 100000_82000_M1 100000_82000_M2 0.050
r 100000_84000_M1 100000_84000_M2 0.050
r 100000_86000_M1 100000_86000_M2 0.050
r 100000_88000_M1 100000_88000_M2 0.050
r 100000_90000_M1 100000_90000_M2 0.050
r 100000_92000_M1 100000_92000_M2 0.050
r 100000_94000_M1 100000_94000_M2 0.050
r 100000_96000_M1 100000_96000_M2 0.050
r 100000_98000_M1 100000_98000_M2 0.050
r 100000_100000_M1 100000_100000_M2 0.050

* ============================================================================
* Via connections M2 to M3
* ============================================================================

r 4000_4000_M2 4000_4000_M3 0.040
r 4000_8000_M2 4000_8000_M3 0.040
r 4000_12000_M2 4000_12000_M3 0.040
r 4000_16000_M2 4000_16000_M3 0.040
r 4000_20000_M2 4000_20000_M3 0.040
r 4000_24000_M2 4000_24000_M3 0.040
r 4000_28000_M2 4000_28000_M3 0.040
r 4000_32000_M2 4000_32000_M3 0.040
r 4000_36000_M2 4000_36000_M3 0.040
r 4000_40000_M2 4000_40000_M3 0.040
r 4000_44000_M2 4000_44000_M3 0.040
r 4000_48000_M2 4000_48000_M3 0.040
r 4000_52000_M2 4000_52000_M3 0.040
r 4000_56000_M2 4000_56000_M3 0.040
r 4000_60000_M2 4000_60000_M3 0.040
r 4000_64000_M2 4000_64000_M3 0.040
r 4000_68000_M2 4000_68000_M3 0.040
r 4000_72000_M2 4000_72000_M3 0.040
r 4000_76000_M2 4000_76000_M3 0.040
r 4000_80000_M2 4000_80000_M3 0.040
r 4000_84000_M2 4000_84000_M3 0.040
r 4000_88000_M2 4000_88000_M3 0.040
r 4000_92000_M2 4000_92000_M3 0.040
r 4000_96000_M2 4000_96000_M3 0.040
r 4000_100000_M2 4000_100000_M3 0.040
r 8000_4000_M2 8000_4000_M3 0.040
r 8000_8000_M2 8000_8000_M3 0.040
r 8000_12000_M2 8000_12000_M3 0.040
r 8000_16000_M2 8000_16000_M3 0.040
r 8000_20000_M2 8000_20000_M3 0.040
r 8000_24000_M2 8000_24000_M3 0.040
r 8000_28000_M2 8000_28000_M3 0.040
r 8000_32000_M2 8000_32000_M3 0.040
r 8000_36000_M2 8000_36000_M3 0.040
r 8000_40000_M2 8000_40000_M3 0.040
r 8000_44000_M2 8000_44000_M3 0.040
r 8000_48000_M2 8000_48000_M3 0.040
r 8000_52000_M2 8000_52000_M3 0.040
r 8000_56000_M2 8000_56000_M3 0.040
r 8000_60000_M2 8000_60000_M3 0.040
r 8000_64000_M2 8000_64000_M3 0.040
r 8000_68000_M2 8000_68000_M3 0.040
r 8000_72000_M2 8000_72000_M3 0.040
r 8000_76000_M2 8000_76000_M3 0.040
r 8000_80000_M2 8000_80000_M3 0.040
r 8000_84000_M2 8000_84000_M3 0.040
r 8000_88000_M2 8000_88000_M3 0.040
r 8000_92000_M2 8000_92000_M3 0.040
r 8000_96000_M2 8000_96000_M3 0.040
r 8000_100000_M2 8000_100000_M3 0.040
r 12000_4000_M2 12000_4000_M3 0.040
r 12000_8000_M2 12000_8000_M3 0.040
r 12000_12000_M2 12000_12000_M3 0.040
r 12000_16000_M2 12000_16000_M3 0.040
r 12000_20000_M2 12000_20000_M3 0.040
r 12000_24000_M2 12000_24000_M3 0.040
r 12000_28000_M2 12000_28000_M3 0.040
r 12000_32000_M2 12000_32000_M3 0.040
r 12000_36000_M2 12000_36000_M3 0.040
r 12000_40000_M2 12000_40000_M3 0.040
r 12000_44000_M2 12000_44000_M3 0.040
r 12000_48000_M2 12000_48000_M3 0.040
r 12000_52000_M2 12000_52000_M3 0.040
r 12000_56000_M2 12000_56000_M3 0.040
r 12000_60000_M2 12000_60000_M3 0.040
r 12000_64000_M2 12000_64000_M3 0.040
r 12000_68000_M2 12000_68000_M3 0.040
r 12000_72000_M2 12000_72000_M3 0.040
r 12000_76000_M2 12000_76000_M3 0.040
r 12000_80000_M2 12000_80000_M3 0.040
r 12000_84000_M2 12000_84000_M3 0.040
r 12000_88000_M2 12000_88000_M3 0.040
r 12000_92000_M2 12000_92000_M3 0.040
r 12000_96000_M2 12000_96000_M3 0.040
r 12000_100000_M2 12000_100000_M3 0.040
r 16000_4000_M2 16000_4000_M3 0.040
r 16000_8000_M2 16000_8000_M3 0.040
r 16000_12000_M2 16000_12000_M3 0.040
r 16000_16000_M2 16000_16000_M3 0.040
r 16000_20000_M2 16000_20000_M3 0.040
r 16000_24000_M2 16000_24000_M3 0.040
r 16000_28000_M2 16000_28000_M3 0.040
r 16000_32000_M2 16000_32000_M3 0.040
r 16000_36000_M2 16000_36000_M3 0.040
r 16000_40000_M2 16000_40000_M3 0.040
r 16000_44000_M2 16000_44000_M3 0.040
r 16000_48000_M2 16000_48000_M3 0.040
r 16000_52000_M2 16000_52000_M3 0.040
r 16000_56000_M2 16000_56000_M3 0.040
r 16000_60000_M2 16000_60000_M3 0.040
r 16000_64000_M2 16000_64000_M3 0.040
r 16000_68000_M2 16000_68000_M3 0.040
r 16000_72000_M2 16000_72000_M3 0.040
r 16000_76000_M2 16000_76000_M3 0.040
r 16000_80000_M2 16000_80000_M3 0.040
r 16000_84000_M2 16000_84000_M3 0.040
r 16000_88000_M2 16000_88000_M3 0.040
r 16000_92000_M2 16000_92000_M3 0.040
r 16000_96000_M2 16000_96000_M3 0.040
r 16000_100000_M2 16000_100000_M3 0.040
r 20000_4000_M2 20000_4000_M3 0.040
r 20000_8000_M2 20000_8000_M3 0.040
r 20000_12000_M2 20000_12000_M3 0.040
r 20000_16000_M2 20000_16000_M3 0.040
r 20000_20000_M2 20000_20000_M3 0.040
r 20000_24000_M2 20000_24000_M3 0.040
r 20000_28000_M2 20000_28000_M3 0.040
r 20000_32000_M2 20000_32000_M3 0.040
r 20000_36000_M2 20000_36000_M3 0.040
r 20000_40000_M2 20000_40000_M3 0.040
r 20000_44000_M2 20000_44000_M3 0.040
r 20000_48000_M2 20000_48000_M3 0.040
r 20000_52000_M2 20000_52000_M3 0.040
r 20000_56000_M2 20000_56000_M3 0.040
r 20000_60000_M2 20000_60000_M3 0.040
r 20000_64000_M2 20000_64000_M3 0.040
r 20000_68000_M2 20000_68000_M3 0.040
r 20000_72000_M2 20000_72000_M3 0.040
r 20000_76000_M2 20000_76000_M3 0.040
r 20000_80000_M2 20000_80000_M3 0.040
r 20000_84000_M2 20000_84000_M3 0.040
r 20000_88000_M2 20000_88000_M3 0.040
r 20000_92000_M2 20000_92000_M3 0.040
r 20000_96000_M2 20000_96000_M3 0.040
r 20000_100000_M2 20000_100000_M3 0.040
r 24000_4000_M2 24000_4000_M3 0.040
r 24000_8000_M2 24000_8000_M3 0.040
r 24000_12000_M2 24000_12000_M3 0.040
r 24000_16000_M2 24000_16000_M3 0.040
r 24000_20000_M2 24000_20000_M3 0.040
r 24000_24000_M2 24000_24000_M3 0.040
r 24000_28000_M2 24000_28000_M3 0.040
r 24000_32000_M2 24000_32000_M3 0.040
r 24000_36000_M2 24000_36000_M3 0.040
r 24000_40000_M2 24000_40000_M3 0.040
r 24000_44000_M2 24000_44000_M3 0.040
r 24000_48000_M2 24000_48000_M3 0.040
r 24000_52000_M2 24000_52000_M3 0.040
r 24000_56000_M2 24000_56000_M3 0.040
r 24000_60000_M2 24000_60000_M3 0.040
r 24000_64000_M2 24000_64000_M3 0.040
r 24000_68000_M2 24000_68000_M3 0.040
r 24000_72000_M2 24000_72000_M3 0.040
r 24000_76000_M2 24000_76000_M3 0.040
r 24000_80000_M2 24000_80000_M3 0.040
r 24000_84000_M2 24000_84000_M3 0.040
r 24000_88000_M2 24000_88000_M3 0.040
r 24000_92000_M2 24000_92000_M3 0.040
r 24000_96000_M2 24000_96000_M3 0.040
r 24000_100000_M2 24000_100000_M3 0.040
r 28000_4000_M2 28000_4000_M3 0.040
r 28000_8000_M2 28000_8000_M3 0.040
r 28000_12000_M2 28000_12000_M3 0.040
r 28000_16000_M2 28000_16000_M3 0.040
r 28000_20000_M2 28000_20000_M3 0.040
r 28000_24000_M2 28000_24000_M3 0.040
r 28000_28000_M2 28000_28000_M3 0.040
r 28000_32000_M2 28000_32000_M3 0.040
r 28000_36000_M2 28000_36000_M3 0.040
r 28000_40000_M2 28000_40000_M3 0.040
r 28000_44000_M2 28000_44000_M3 0.040
r 28000_48000_M2 28000_48000_M3 0.040
r 28000_52000_M2 28000_52000_M3 0.040
r 28000_56000_M2 28000_56000_M3 0.040
r 28000_60000_M2 28000_60000_M3 0.040
r 28000_64000_M2 28000_64000_M3 0.040
r 28000_68000_M2 28000_68000_M3 0.040
r 28000_72000_M2 28000_72000_M3 0.040
r 28000_76000_M2 28000_76000_M3 0.040
r 28000_80000_M2 28000_80000_M3 0.040
r 28000_84000_M2 28000_84000_M3 0.040
r 28000_88000_M2 28000_88000_M3 0.040
r 28000_92000_M2 28000_92000_M3 0.040
r 28000_96000_M2 28000_96000_M3 0.040
r 28000_100000_M2 28000_100000_M3 0.040
r 32000_4000_M2 32000_4000_M3 0.040
r 32000_8000_M2 32000_8000_M3 0.040
r 32000_12000_M2 32000_12000_M3 0.040
r 32000_16000_M2 32000_16000_M3 0.040
r 32000_20000_M2 32000_20000_M3 0.040
r 32000_24000_M2 32000_24000_M3 0.040
r 32000_28000_M2 32000_28000_M3 0.040
r 32000_32000_M2 32000_32000_M3 0.040
r 32000_36000_M2 32000_36000_M3 0.040
r 32000_40000_M2 32000_40000_M3 0.040
r 32000_44000_M2 32000_44000_M3 0.040
r 32000_48000_M2 32000_48000_M3 0.040
r 32000_52000_M2 32000_52000_M3 0.040
r 32000_56000_M2 32000_56000_M3 0.040
r 32000_60000_M2 32000_60000_M3 0.040
r 32000_64000_M2 32000_64000_M3 0.040
r 32000_68000_M2 32000_68000_M3 0.040
r 32000_72000_M2 32000_72000_M3 0.040
r 32000_76000_M2 32000_76000_M3 0.040
r 32000_80000_M2 32000_80000_M3 0.040
r 32000_84000_M2 32000_84000_M3 0.040
r 32000_88000_M2 32000_88000_M3 0.040
r 32000_92000_M2 32000_92000_M3 0.040
r 32000_96000_M2 32000_96000_M3 0.040
r 32000_100000_M2 32000_100000_M3 0.040
r 36000_4000_M2 36000_4000_M3 0.040
r 36000_8000_M2 36000_8000_M3 0.040
r 36000_12000_M2 36000_12000_M3 0.040
r 36000_16000_M2 36000_16000_M3 0.040
r 36000_20000_M2 36000_20000_M3 0.040
r 36000_24000_M2 36000_24000_M3 0.040
r 36000_28000_M2 36000_28000_M3 0.040
r 36000_32000_M2 36000_32000_M3 0.040
r 36000_36000_M2 36000_36000_M3 0.040
r 36000_40000_M2 36000_40000_M3 0.040
r 36000_44000_M2 36000_44000_M3 0.040
r 36000_48000_M2 36000_48000_M3 0.040
r 36000_52000_M2 36000_52000_M3 0.040
r 36000_56000_M2 36000_56000_M3 0.040
r 36000_60000_M2 36000_60000_M3 0.040
r 36000_64000_M2 36000_64000_M3 0.040
r 36000_68000_M2 36000_68000_M3 0.040
r 36000_72000_M2 36000_72000_M3 0.040
r 36000_76000_M2 36000_76000_M3 0.040
r 36000_80000_M2 36000_80000_M3 0.040
r 36000_84000_M2 36000_84000_M3 0.040
r 36000_88000_M2 36000_88000_M3 0.040
r 36000_92000_M2 36000_92000_M3 0.040
r 36000_96000_M2 36000_96000_M3 0.040
r 36000_100000_M2 36000_100000_M3 0.040
r 40000_4000_M2 40000_4000_M3 0.040
r 40000_8000_M2 40000_8000_M3 0.040
r 40000_12000_M2 40000_12000_M3 0.040
r 40000_16000_M2 40000_16000_M3 0.040
r 40000_20000_M2 40000_20000_M3 0.040
r 40000_24000_M2 40000_24000_M3 0.040
r 40000_28000_M2 40000_28000_M3 0.040
r 40000_32000_M2 40000_32000_M3 0.040
r 40000_36000_M2 40000_36000_M3 0.040
r 40000_40000_M2 40000_40000_M3 0.040
r 40000_44000_M2 40000_44000_M3 0.040
r 40000_48000_M2 40000_48000_M3 0.040
r 40000_52000_M2 40000_52000_M3 0.040
r 40000_56000_M2 40000_56000_M3 0.040
r 40000_60000_M2 40000_60000_M3 0.040
r 40000_64000_M2 40000_64000_M3 0.040
r 40000_68000_M2 40000_68000_M3 0.040
r 40000_72000_M2 40000_72000_M3 0.040
r 40000_76000_M2 40000_76000_M3 0.040
r 40000_80000_M2 40000_80000_M3 0.040
r 40000_84000_M2 40000_84000_M3 0.040
r 40000_88000_M2 40000_88000_M3 0.040
r 40000_92000_M2 40000_92000_M3 0.040
r 40000_96000_M2 40000_96000_M3 0.040
r 40000_100000_M2 40000_100000_M3 0.040
r 44000_4000_M2 44000_4000_M3 0.040
r 44000_8000_M2 44000_8000_M3 0.040
r 44000_12000_M2 44000_12000_M3 0.040
r 44000_16000_M2 44000_16000_M3 0.040
r 44000_20000_M2 44000_20000_M3 0.040
r 44000_24000_M2 44000_24000_M3 0.040
r 44000_28000_M2 44000_28000_M3 0.040
r 44000_32000_M2 44000_32000_M3 0.040
r 44000_36000_M2 44000_36000_M3 0.040
r 44000_40000_M2 44000_40000_M3 0.040
r 44000_44000_M2 44000_44000_M3 0.040
r 44000_48000_M2 44000_48000_M3 0.040
r 44000_52000_M2 44000_52000_M3 0.040
r 44000_56000_M2 44000_56000_M3 0.040
r 44000_60000_M2 44000_60000_M3 0.040
r 44000_64000_M2 44000_64000_M3 0.040
r 44000_68000_M2 44000_68000_M3 0.040
r 44000_72000_M2 44000_72000_M3 0.040
r 44000_76000_M2 44000_76000_M3 0.040
r 44000_80000_M2 44000_80000_M3 0.040
r 44000_84000_M2 44000_84000_M3 0.040
r 44000_88000_M2 44000_88000_M3 0.040
r 44000_92000_M2 44000_92000_M3 0.040
r 44000_96000_M2 44000_96000_M3 0.040
r 44000_100000_M2 44000_100000_M3 0.040
r 48000_4000_M2 48000_4000_M3 0.040
r 48000_8000_M2 48000_8000_M3 0.040
r 48000_12000_M2 48000_12000_M3 0.040
r 48000_16000_M2 48000_16000_M3 0.040
r 48000_20000_M2 48000_20000_M3 0.040
r 48000_24000_M2 48000_24000_M3 0.040
r 48000_28000_M2 48000_28000_M3 0.040
r 48000_32000_M2 48000_32000_M3 0.040
r 48000_36000_M2 48000_36000_M3 0.040
r 48000_40000_M2 48000_40000_M3 0.040
r 48000_44000_M2 48000_44000_M3 0.040
r 48000_48000_M2 48000_48000_M3 0.040
r 48000_52000_M2 48000_52000_M3 0.040
r 48000_56000_M2 48000_56000_M3 0.040
r 48000_60000_M2 48000_60000_M3 0.040
r 48000_64000_M2 48000_64000_M3 0.040
r 48000_68000_M2 48000_68000_M3 0.040
r 48000_72000_M2 48000_72000_M3 0.040
r 48000_76000_M2 48000_76000_M3 0.040
r 48000_80000_M2 48000_80000_M3 0.040
r 48000_84000_M2 48000_84000_M3 0.040
r 48000_88000_M2 48000_88000_M3 0.040
r 48000_92000_M2 48000_92000_M3 0.040
r 48000_96000_M2 48000_96000_M3 0.040
r 48000_100000_M2 48000_100000_M3 0.040
r 52000_4000_M2 52000_4000_M3 0.040
r 52000_8000_M2 52000_8000_M3 0.040
r 52000_12000_M2 52000_12000_M3 0.040
r 52000_16000_M2 52000_16000_M3 0.040
r 52000_20000_M2 52000_20000_M3 0.040
r 52000_24000_M2 52000_24000_M3 0.040
r 52000_28000_M2 52000_28000_M3 0.040
r 52000_32000_M2 52000_32000_M3 0.040
r 52000_36000_M2 52000_36000_M3 0.040
r 52000_40000_M2 52000_40000_M3 0.040
r 52000_44000_M2 52000_44000_M3 0.040
r 52000_48000_M2 52000_48000_M3 0.040
r 52000_52000_M2 52000_52000_M3 0.040
r 52000_56000_M2 52000_56000_M3 0.040
r 52000_60000_M2 52000_60000_M3 0.040
r 52000_64000_M2 52000_64000_M3 0.040
r 52000_68000_M2 52000_68000_M3 0.040
r 52000_72000_M2 52000_72000_M3 0.040
r 52000_76000_M2 52000_76000_M3 0.040
r 52000_80000_M2 52000_80000_M3 0.040
r 52000_84000_M2 52000_84000_M3 0.040
r 52000_88000_M2 52000_88000_M3 0.040
r 52000_92000_M2 52000_92000_M3 0.040
r 52000_96000_M2 52000_96000_M3 0.040
r 52000_100000_M2 52000_100000_M3 0.040
r 56000_4000_M2 56000_4000_M3 0.040
r 56000_8000_M2 56000_8000_M3 0.040
r 56000_12000_M2 56000_12000_M3 0.040
r 56000_16000_M2 56000_16000_M3 0.040
r 56000_20000_M2 56000_20000_M3 0.040
r 56000_24000_M2 56000_24000_M3 0.040
r 56000_28000_M2 56000_28000_M3 0.040
r 56000_32000_M2 56000_32000_M3 0.040
r 56000_36000_M2 56000_36000_M3 0.040
r 56000_40000_M2 56000_40000_M3 0.040
r 56000_44000_M2 56000_44000_M3 0.040
r 56000_48000_M2 56000_48000_M3 0.040
r 56000_52000_M2 56000_52000_M3 0.040
r 56000_56000_M2 56000_56000_M3 0.040
r 56000_60000_M2 56000_60000_M3 0.040
r 56000_64000_M2 56000_64000_M3 0.040
r 56000_68000_M2 56000_68000_M3 0.040
r 56000_72000_M2 56000_72000_M3 0.040
r 56000_76000_M2 56000_76000_M3 0.040
r 56000_80000_M2 56000_80000_M3 0.040
r 56000_84000_M2 56000_84000_M3 0.040
r 56000_88000_M2 56000_88000_M3 0.040
r 56000_92000_M2 56000_92000_M3 0.040
r 56000_96000_M2 56000_96000_M3 0.040
r 56000_100000_M2 56000_100000_M3 0.040
r 60000_4000_M2 60000_4000_M3 0.040
r 60000_8000_M2 60000_8000_M3 0.040
r 60000_12000_M2 60000_12000_M3 0.040
r 60000_16000_M2 60000_16000_M3 0.040
r 60000_20000_M2 60000_20000_M3 0.040
r 60000_24000_M2 60000_24000_M3 0.040
r 60000_28000_M2 60000_28000_M3 0.040
r 60000_32000_M2 60000_32000_M3 0.040
r 60000_36000_M2 60000_36000_M3 0.040
r 60000_40000_M2 60000_40000_M3 0.040
r 60000_44000_M2 60000_44000_M3 0.040
r 60000_48000_M2 60000_48000_M3 0.040
r 60000_52000_M2 60000_52000_M3 0.040
r 60000_56000_M2 60000_56000_M3 0.040
r 60000_60000_M2 60000_60000_M3 0.040
r 60000_64000_M2 60000_64000_M3 0.040
r 60000_68000_M2 60000_68000_M3 0.040
r 60000_72000_M2 60000_72000_M3 0.040
r 60000_76000_M2 60000_76000_M3 0.040
r 60000_80000_M2 60000_80000_M3 0.040
r 60000_84000_M2 60000_84000_M3 0.040
r 60000_88000_M2 60000_88000_M3 0.040
r 60000_92000_M2 60000_92000_M3 0.040
r 60000_96000_M2 60000_96000_M3 0.040
r 60000_100000_M2 60000_100000_M3 0.040
r 64000_4000_M2 64000_4000_M3 0.040
r 64000_8000_M2 64000_8000_M3 0.040
r 64000_12000_M2 64000_12000_M3 0.040
r 64000_16000_M2 64000_16000_M3 0.040
r 64000_20000_M2 64000_20000_M3 0.040
r 64000_24000_M2 64000_24000_M3 0.040
r 64000_28000_M2 64000_28000_M3 0.040
r 64000_32000_M2 64000_32000_M3 0.040
r 64000_36000_M2 64000_36000_M3 0.040
r 64000_40000_M2 64000_40000_M3 0.040
r 64000_44000_M2 64000_44000_M3 0.040
r 64000_48000_M2 64000_48000_M3 0.040
r 64000_52000_M2 64000_52000_M3 0.040
r 64000_56000_M2 64000_56000_M3 0.040
r 64000_60000_M2 64000_60000_M3 0.040
r 64000_64000_M2 64000_64000_M3 0.040
r 64000_68000_M2 64000_68000_M3 0.040
r 64000_72000_M2 64000_72000_M3 0.040
r 64000_76000_M2 64000_76000_M3 0.040
r 64000_80000_M2 64000_80000_M3 0.040
r 64000_84000_M2 64000_84000_M3 0.040
r 64000_88000_M2 64000_88000_M3 0.040
r 64000_92000_M2 64000_92000_M3 0.040
r 64000_96000_M2 64000_96000_M3 0.040
r 64000_100000_M2 64000_100000_M3 0.040
r 68000_4000_M2 68000_4000_M3 0.040
r 68000_8000_M2 68000_8000_M3 0.040
r 68000_12000_M2 68000_12000_M3 0.040
r 68000_16000_M2 68000_16000_M3 0.040
r 68000_20000_M2 68000_20000_M3 0.040
r 68000_24000_M2 68000_24000_M3 0.040
r 68000_28000_M2 68000_28000_M3 0.040
r 68000_32000_M2 68000_32000_M3 0.040
r 68000_36000_M2 68000_36000_M3 0.040
r 68000_40000_M2 68000_40000_M3 0.040
r 68000_44000_M2 68000_44000_M3 0.040
r 68000_48000_M2 68000_48000_M3 0.040
r 68000_52000_M2 68000_52000_M3 0.040
r 68000_56000_M2 68000_56000_M3 0.040
r 68000_60000_M2 68000_60000_M3 0.040
r 68000_64000_M2 68000_64000_M3 0.040
r 68000_68000_M2 68000_68000_M3 0.040
r 68000_72000_M2 68000_72000_M3 0.040
r 68000_76000_M2 68000_76000_M3 0.040
r 68000_80000_M2 68000_80000_M3 0.040
r 68000_84000_M2 68000_84000_M3 0.040
r 68000_88000_M2 68000_88000_M3 0.040
r 68000_92000_M2 68000_92000_M3 0.040
r 68000_96000_M2 68000_96000_M3 0.040
r 68000_100000_M2 68000_100000_M3 0.040
r 72000_4000_M2 72000_4000_M3 0.040
r 72000_8000_M2 72000_8000_M3 0.040
r 72000_12000_M2 72000_12000_M3 0.040
r 72000_16000_M2 72000_16000_M3 0.040
r 72000_20000_M2 72000_20000_M3 0.040
r 72000_24000_M2 72000_24000_M3 0.040
r 72000_28000_M2 72000_28000_M3 0.040
r 72000_32000_M2 72000_32000_M3 0.040
r 72000_36000_M2 72000_36000_M3 0.040
r 72000_40000_M2 72000_40000_M3 0.040
r 72000_44000_M2 72000_44000_M3 0.040
r 72000_48000_M2 72000_48000_M3 0.040
r 72000_52000_M2 72000_52000_M3 0.040
r 72000_56000_M2 72000_56000_M3 0.040
r 72000_60000_M2 72000_60000_M3 0.040
r 72000_64000_M2 72000_64000_M3 0.040
r 72000_68000_M2 72000_68000_M3 0.040
r 72000_72000_M2 72000_72000_M3 0.040
r 72000_76000_M2 72000_76000_M3 0.040
r 72000_80000_M2 72000_80000_M3 0.040
r 72000_84000_M2 72000_84000_M3 0.040
r 72000_88000_M2 72000_88000_M3 0.040
r 72000_92000_M2 72000_92000_M3 0.040
r 72000_96000_M2 72000_96000_M3 0.040
r 72000_100000_M2 72000_100000_M3 0.040
r 76000_4000_M2 76000_4000_M3 0.040
r 76000_8000_M2 76000_8000_M3 0.040
r 76000_12000_M2 76000_12000_M3 0.040
r 76000_16000_M2 76000_16000_M3 0.040
r 76000_20000_M2 76000_20000_M3 0.040
r 76000_24000_M2 76000_24000_M3 0.040
r 76000_28000_M2 76000_28000_M3 0.040
r 76000_32000_M2 76000_32000_M3 0.040
r 76000_36000_M2 76000_36000_M3 0.040
r 76000_40000_M2 76000_40000_M3 0.040
r 76000_44000_M2 76000_44000_M3 0.040
r 76000_48000_M2 76000_48000_M3 0.040
r 76000_52000_M2 76000_52000_M3 0.040
r 76000_56000_M2 76000_56000_M3 0.040
r 76000_60000_M2 76000_60000_M3 0.040
r 76000_64000_M2 76000_64000_M3 0.040
r 76000_68000_M2 76000_68000_M3 0.040
r 76000_72000_M2 76000_72000_M3 0.040
r 76000_76000_M2 76000_76000_M3 0.040
r 76000_80000_M2 76000_80000_M3 0.040
r 76000_84000_M2 76000_84000_M3 0.040
r 76000_88000_M2 76000_88000_M3 0.040
r 76000_92000_M2 76000_92000_M3 0.040
r 76000_96000_M2 76000_96000_M3 0.040
r 76000_100000_M2 76000_100000_M3 0.040
r 80000_4000_M2 80000_4000_M3 0.040
r 80000_8000_M2 80000_8000_M3 0.040
r 80000_12000_M2 80000_12000_M3 0.040
r 80000_16000_M2 80000_16000_M3 0.040
r 80000_20000_M2 80000_20000_M3 0.040
r 80000_24000_M2 80000_24000_M3 0.040
r 80000_28000_M2 80000_28000_M3 0.040
r 80000_32000_M2 80000_32000_M3 0.040
r 80000_36000_M2 80000_36000_M3 0.040
r 80000_40000_M2 80000_40000_M3 0.040
r 80000_44000_M2 80000_44000_M3 0.040
r 80000_48000_M2 80000_48000_M3 0.040
r 80000_52000_M2 80000_52000_M3 0.040
r 80000_56000_M2 80000_56000_M3 0.040
r 80000_60000_M2 80000_60000_M3 0.040
r 80000_64000_M2 80000_64000_M3 0.040
r 80000_68000_M2 80000_68000_M3 0.040
r 80000_72000_M2 80000_72000_M3 0.040
r 80000_76000_M2 80000_76000_M3 0.040
r 80000_80000_M2 80000_80000_M3 0.040
r 80000_84000_M2 80000_84000_M3 0.040
r 80000_88000_M2 80000_88000_M3 0.040
r 80000_92000_M2 80000_92000_M3 0.040
r 80000_96000_M2 80000_96000_M3 0.040
r 80000_100000_M2 80000_100000_M3 0.040
r 84000_4000_M2 84000_4000_M3 0.040
r 84000_8000_M2 84000_8000_M3 0.040
r 84000_12000_M2 84000_12000_M3 0.040
r 84000_16000_M2 84000_16000_M3 0.040
r 84000_20000_M2 84000_20000_M3 0.040
r 84000_24000_M2 84000_24000_M3 0.040
r 84000_28000_M2 84000_28000_M3 0.040
r 84000_32000_M2 84000_32000_M3 0.040
r 84000_36000_M2 84000_36000_M3 0.040
r 84000_40000_M2 84000_40000_M3 0.040
r 84000_44000_M2 84000_44000_M3 0.040
r 84000_48000_M2 84000_48000_M3 0.040
r 84000_52000_M2 84000_52000_M3 0.040
r 84000_56000_M2 84000_56000_M3 0.040
r 84000_60000_M2 84000_60000_M3 0.040
r 84000_64000_M2 84000_64000_M3 0.040
r 84000_68000_M2 84000_68000_M3 0.040
r 84000_72000_M2 84000_72000_M3 0.040
r 84000_76000_M2 84000_76000_M3 0.040
r 84000_80000_M2 84000_80000_M3 0.040
r 84000_84000_M2 84000_84000_M3 0.040
r 84000_88000_M2 84000_88000_M3 0.040
r 84000_92000_M2 84000_92000_M3 0.040
r 84000_96000_M2 84000_96000_M3 0.040
r 84000_100000_M2 84000_100000_M3 0.040
r 88000_4000_M2 88000_4000_M3 0.040
r 88000_8000_M2 88000_8000_M3 0.040
r 88000_12000_M2 88000_12000_M3 0.040
r 88000_16000_M2 88000_16000_M3 0.040
r 88000_20000_M2 88000_20000_M3 0.040
r 88000_24000_M2 88000_24000_M3 0.040
r 88000_28000_M2 88000_28000_M3 0.040
r 88000_32000_M2 88000_32000_M3 0.040
r 88000_36000_M2 88000_36000_M3 0.040
r 88000_40000_M2 88000_40000_M3 0.040
r 88000_44000_M2 88000_44000_M3 0.040
r 88000_48000_M2 88000_48000_M3 0.040
r 88000_52000_M2 88000_52000_M3 0.040
r 88000_56000_M2 88000_56000_M3 0.040
r 88000_60000_M2 88000_60000_M3 0.040
r 88000_64000_M2 88000_64000_M3 0.040
r 88000_68000_M2 88000_68000_M3 0.040
r 88000_72000_M2 88000_72000_M3 0.040
r 88000_76000_M2 88000_76000_M3 0.040
r 88000_80000_M2 88000_80000_M3 0.040
r 88000_84000_M2 88000_84000_M3 0.040
r 88000_88000_M2 88000_88000_M3 0.040
r 88000_92000_M2 88000_92000_M3 0.040
r 88000_96000_M2 88000_96000_M3 0.040
r 88000_100000_M2 88000_100000_M3 0.040
r 92000_4000_M2 92000_4000_M3 0.040
r 92000_8000_M2 92000_8000_M3 0.040
r 92000_12000_M2 92000_12000_M3 0.040
r 92000_16000_M2 92000_16000_M3 0.040
r 92000_20000_M2 92000_20000_M3 0.040
r 92000_24000_M2 92000_24000_M3 0.040
r 92000_28000_M2 92000_28000_M3 0.040
r 92000_32000_M2 92000_32000_M3 0.040
r 92000_36000_M2 92000_36000_M3 0.040
r 92000_40000_M2 92000_40000_M3 0.040
r 92000_44000_M2 92000_44000_M3 0.040
r 92000_48000_M2 92000_48000_M3 0.040
r 92000_52000_M2 92000_52000_M3 0.040
r 92000_56000_M2 92000_56000_M3 0.040
r 92000_60000_M2 92000_60000_M3 0.040
r 92000_64000_M2 92000_64000_M3 0.040
r 92000_68000_M2 92000_68000_M3 0.040
r 92000_72000_M2 92000_72000_M3 0.040
r 92000_76000_M2 92000_76000_M3 0.040
r 92000_80000_M2 92000_80000_M3 0.040
r 92000_84000_M2 92000_84000_M3 0.040
r 92000_88000_M2 92000_88000_M3 0.040
r 92000_92000_M2 92000_92000_M3 0.040
r 92000_96000_M2 92000_96000_M3 0.040
r 92000_100000_M2 92000_100000_M3 0.040
r 96000_4000_M2 96000_4000_M3 0.040
r 96000_8000_M2 96000_8000_M3 0.040
r 96000_12000_M2 96000_12000_M3 0.040
r 96000_16000_M2 96000_16000_M3 0.040
r 96000_20000_M2 96000_20000_M3 0.040
r 96000_24000_M2 96000_24000_M3 0.040
r 96000_28000_M2 96000_28000_M3 0.040
r 96000_32000_M2 96000_32000_M3 0.040
r 96000_36000_M2 96000_36000_M3 0.040
r 96000_40000_M2 96000_40000_M3 0.040
r 96000_44000_M2 96000_44000_M3 0.040
r 96000_48000_M2 96000_48000_M3 0.040
r 96000_52000_M2 96000_52000_M3 0.040
r 96000_56000_M2 96000_56000_M3 0.040
r 96000_60000_M2 96000_60000_M3 0.040
r 96000_64000_M2 96000_64000_M3 0.040
r 96000_68000_M2 96000_68000_M3 0.040
r 96000_72000_M2 96000_72000_M3 0.040
r 96000_76000_M2 96000_76000_M3 0.040
r 96000_80000_M2 96000_80000_M3 0.040
r 96000_84000_M2 96000_84000_M3 0.040
r 96000_88000_M2 96000_88000_M3 0.040
r 96000_92000_M2 96000_92000_M3 0.040
r 96000_96000_M2 96000_96000_M3 0.040
r 96000_100000_M2 96000_100000_M3 0.040
r 100000_4000_M2 100000_4000_M3 0.040
r 100000_8000_M2 100000_8000_M3 0.040
r 100000_12000_M2 100000_12000_M3 0.040
r 100000_16000_M2 100000_16000_M3 0.040
r 100000_20000_M2 100000_20000_M3 0.040
r 100000_24000_M2 100000_24000_M3 0.040
r 100000_28000_M2 100000_28000_M3 0.040
r 100000_32000_M2 100000_32000_M3 0.040
r 100000_36000_M2 100000_36000_M3 0.040
r 100000_40000_M2 100000_40000_M3 0.040
r 100000_44000_M2 100000_44000_M3 0.040
r 100000_48000_M2 100000_48000_M3 0.040
r 100000_52000_M2 100000_52000_M3 0.040
r 100000_56000_M2 100000_56000_M3 0.040
r 100000_60000_M2 100000_60000_M3 0.040
r 100000_64000_M2 100000_64000_M3 0.040
r 100000_68000_M2 100000_68000_M3 0.040
r 100000_72000_M2 100000_72000_M3 0.040
r 100000_76000_M2 100000_76000_M3 0.040
r 100000_80000_M2 100000_80000_M3 0.040
r 100000_84000_M2 100000_84000_M3 0.040
r 100000_88000_M2 100000_88000_M3 0.040
r 100000_92000_M2 100000_92000_M3 0.040
r 100000_96000_M2 100000_96000_M3 0.040
r 100000_100000_M2 100000_100000_M3 0.040

* ============================================================================
* Via connections M3 to M4
* ============================================================================

r 4000_4000_M3 4000_4000_M4 0.035
r 4000_8000_M3 4000_8000_M4 0.035
r 4000_12000_M3 4000_12000_M4 0.035
r 4000_16000_M3 4000_16000_M4 0.035
r 4000_20000_M3 4000_20000_M4 0.035
r 4000_24000_M3 4000_24000_M4 0.035
r 4000_28000_M3 4000_28000_M4 0.035
r 4000_32000_M3 4000_32000_M4 0.035
r 4000_36000_M3 4000_36000_M4 0.035
r 4000_40000_M3 4000_40000_M4 0.035
r 4000_44000_M3 4000_44000_M4 0.035
r 4000_48000_M3 4000_48000_M4 0.035
r 4000_52000_M3 4000_52000_M4 0.035
r 4000_56000_M3 4000_56000_M4 0.035
r 4000_60000_M3 4000_60000_M4 0.035
r 4000_64000_M3 4000_64000_M4 0.035
r 4000_68000_M3 4000_68000_M4 0.035
r 4000_72000_M3 4000_72000_M4 0.035
r 4000_76000_M3 4000_76000_M4 0.035
r 4000_80000_M3 4000_80000_M4 0.035
r 4000_84000_M3 4000_84000_M4 0.035
r 4000_88000_M3 4000_88000_M4 0.035
r 4000_92000_M3 4000_92000_M4 0.035
r 4000_96000_M3 4000_96000_M4 0.035
r 4000_100000_M3 4000_100000_M4 0.035
r 8000_4000_M3 8000_4000_M4 0.035
r 8000_8000_M3 8000_8000_M4 0.035
r 8000_12000_M3 8000_12000_M4 0.035
r 8000_16000_M3 8000_16000_M4 0.035
r 8000_20000_M3 8000_20000_M4 0.035
r 8000_24000_M3 8000_24000_M4 0.035
r 8000_28000_M3 8000_28000_M4 0.035
r 8000_32000_M3 8000_32000_M4 0.035
r 8000_36000_M3 8000_36000_M4 0.035
r 8000_40000_M3 8000_40000_M4 0.035
r 8000_44000_M3 8000_44000_M4 0.035
r 8000_48000_M3 8000_48000_M4 0.035
r 8000_52000_M3 8000_52000_M4 0.035
r 8000_56000_M3 8000_56000_M4 0.035
r 8000_60000_M3 8000_60000_M4 0.035
r 8000_64000_M3 8000_64000_M4 0.035
r 8000_68000_M3 8000_68000_M4 0.035
r 8000_72000_M3 8000_72000_M4 0.035
r 8000_76000_M3 8000_76000_M4 0.035
r 8000_80000_M3 8000_80000_M4 0.035
r 8000_84000_M3 8000_84000_M4 0.035
r 8000_88000_M3 8000_88000_M4 0.035
r 8000_92000_M3 8000_92000_M4 0.035
r 8000_96000_M3 8000_96000_M4 0.035
r 8000_100000_M3 8000_100000_M4 0.035
r 12000_4000_M3 12000_4000_M4 0.035
r 12000_8000_M3 12000_8000_M4 0.035
r 12000_12000_M3 12000_12000_M4 0.035
r 12000_16000_M3 12000_16000_M4 0.035
r 12000_20000_M3 12000_20000_M4 0.035
r 12000_24000_M3 12000_24000_M4 0.035
r 12000_28000_M3 12000_28000_M4 0.035
r 12000_32000_M3 12000_32000_M4 0.035
r 12000_36000_M3 12000_36000_M4 0.035
r 12000_40000_M3 12000_40000_M4 0.035
r 12000_44000_M3 12000_44000_M4 0.035
r 12000_48000_M3 12000_48000_M4 0.035
r 12000_52000_M3 12000_52000_M4 0.035
r 12000_56000_M3 12000_56000_M4 0.035
r 12000_60000_M3 12000_60000_M4 0.035
r 12000_64000_M3 12000_64000_M4 0.035
r 12000_68000_M3 12000_68000_M4 0.035
r 12000_72000_M3 12000_72000_M4 0.035
r 12000_76000_M3 12000_76000_M4 0.035
r 12000_80000_M3 12000_80000_M4 0.035
r 12000_84000_M3 12000_84000_M4 0.035
r 12000_88000_M3 12000_88000_M4 0.035
r 12000_92000_M3 12000_92000_M4 0.035
r 12000_96000_M3 12000_96000_M4 0.035
r 12000_100000_M3 12000_100000_M4 0.035
r 16000_4000_M3 16000_4000_M4 0.035
r 16000_8000_M3 16000_8000_M4 0.035
r 16000_12000_M3 16000_12000_M4 0.035
r 16000_16000_M3 16000_16000_M4 0.035
r 16000_20000_M3 16000_20000_M4 0.035
r 16000_24000_M3 16000_24000_M4 0.035
r 16000_28000_M3 16000_28000_M4 0.035
r 16000_32000_M3 16000_32000_M4 0.035
r 16000_36000_M3 16000_36000_M4 0.035
r 16000_40000_M3 16000_40000_M4 0.035
r 16000_44000_M3 16000_44000_M4 0.035
r 16000_48000_M3 16000_48000_M4 0.035
r 16000_52000_M3 16000_52000_M4 0.035
r 16000_56000_M3 16000_56000_M4 0.035
r 16000_60000_M3 16000_60000_M4 0.035
r 16000_64000_M3 16000_64000_M4 0.035
r 16000_68000_M3 16000_68000_M4 0.035
r 16000_72000_M3 16000_72000_M4 0.035
r 16000_76000_M3 16000_76000_M4 0.035
r 16000_80000_M3 16000_80000_M4 0.035
r 16000_84000_M3 16000_84000_M4 0.035
r 16000_88000_M3 16000_88000_M4 0.035
r 16000_92000_M3 16000_92000_M4 0.035
r 16000_96000_M3 16000_96000_M4 0.035
r 16000_100000_M3 16000_100000_M4 0.035
r 20000_4000_M3 20000_4000_M4 0.035
r 20000_8000_M3 20000_8000_M4 0.035
r 20000_12000_M3 20000_12000_M4 0.035
r 20000_16000_M3 20000_16000_M4 0.035
r 20000_20000_M3 20000_20000_M4 0.035
r 20000_24000_M3 20000_24000_M4 0.035
r 20000_28000_M3 20000_28000_M4 0.035
r 20000_32000_M3 20000_32000_M4 0.035
r 20000_36000_M3 20000_36000_M4 0.035
r 20000_40000_M3 20000_40000_M4 0.035
r 20000_44000_M3 20000_44000_M4 0.035
r 20000_48000_M3 20000_48000_M4 0.035
r 20000_52000_M3 20000_52000_M4 0.035
r 20000_56000_M3 20000_56000_M4 0.035
r 20000_60000_M3 20000_60000_M4 0.035
r 20000_64000_M3 20000_64000_M4 0.035
r 20000_68000_M3 20000_68000_M4 0.035
r 20000_72000_M3 20000_72000_M4 0.035
r 20000_76000_M3 20000_76000_M4 0.035
r 20000_80000_M3 20000_80000_M4 0.035
r 20000_84000_M3 20000_84000_M4 0.035
r 20000_88000_M3 20000_88000_M4 0.035
r 20000_92000_M3 20000_92000_M4 0.035
r 20000_96000_M3 20000_96000_M4 0.035
r 20000_100000_M3 20000_100000_M4 0.035
r 24000_4000_M3 24000_4000_M4 0.035
r 24000_8000_M3 24000_8000_M4 0.035
r 24000_12000_M3 24000_12000_M4 0.035
r 24000_16000_M3 24000_16000_M4 0.035
r 24000_20000_M3 24000_20000_M4 0.035
r 24000_24000_M3 24000_24000_M4 0.035
r 24000_28000_M3 24000_28000_M4 0.035
r 24000_32000_M3 24000_32000_M4 0.035
r 24000_36000_M3 24000_36000_M4 0.035
r 24000_40000_M3 24000_40000_M4 0.035
r 24000_44000_M3 24000_44000_M4 0.035
r 24000_48000_M3 24000_48000_M4 0.035
r 24000_52000_M3 24000_52000_M4 0.035
r 24000_56000_M3 24000_56000_M4 0.035
r 24000_60000_M3 24000_60000_M4 0.035
r 24000_64000_M3 24000_64000_M4 0.035
r 24000_68000_M3 24000_68000_M4 0.035
r 24000_72000_M3 24000_72000_M4 0.035
r 24000_76000_M3 24000_76000_M4 0.035
r 24000_80000_M3 24000_80000_M4 0.035
r 24000_84000_M3 24000_84000_M4 0.035
r 24000_88000_M3 24000_88000_M4 0.035
r 24000_92000_M3 24000_92000_M4 0.035
r 24000_96000_M3 24000_96000_M4 0.035
r 24000_100000_M3 24000_100000_M4 0.035
r 28000_4000_M3 28000_4000_M4 0.035
r 28000_8000_M3 28000_8000_M4 0.035
r 28000_12000_M3 28000_12000_M4 0.035
r 28000_16000_M3 28000_16000_M4 0.035
r 28000_20000_M3 28000_20000_M4 0.035
r 28000_24000_M3 28000_24000_M4 0.035
r 28000_28000_M3 28000_28000_M4 0.035
r 28000_32000_M3 28000_32000_M4 0.035
r 28000_36000_M3 28000_36000_M4 0.035
r 28000_40000_M3 28000_40000_M4 0.035
r 28000_44000_M3 28000_44000_M4 0.035
r 28000_48000_M3 28000_48000_M4 0.035
r 28000_52000_M3 28000_52000_M4 0.035
r 28000_56000_M3 28000_56000_M4 0.035
r 28000_60000_M3 28000_60000_M4 0.035
r 28000_64000_M3 28000_64000_M4 0.035
r 28000_68000_M3 28000_68000_M4 0.035
r 28000_72000_M3 28000_72000_M4 0.035
r 28000_76000_M3 28000_76000_M4 0.035
r 28000_80000_M3 28000_80000_M4 0.035
r 28000_84000_M3 28000_84000_M4 0.035
r 28000_88000_M3 28000_88000_M4 0.035
r 28000_92000_M3 28000_92000_M4 0.035
r 28000_96000_M3 28000_96000_M4 0.035
r 28000_100000_M3 28000_100000_M4 0.035
r 32000_4000_M3 32000_4000_M4 0.035
r 32000_8000_M3 32000_8000_M4 0.035
r 32000_12000_M3 32000_12000_M4 0.035
r 32000_16000_M3 32000_16000_M4 0.035
r 32000_20000_M3 32000_20000_M4 0.035
r 32000_24000_M3 32000_24000_M4 0.035
r 32000_28000_M3 32000_28000_M4 0.035
r 32000_32000_M3 32000_32000_M4 0.035
r 32000_36000_M3 32000_36000_M4 0.035
r 32000_40000_M3 32000_40000_M4 0.035
r 32000_44000_M3 32000_44000_M4 0.035
r 32000_48000_M3 32000_48000_M4 0.035
r 32000_52000_M3 32000_52000_M4 0.035
r 32000_56000_M3 32000_56000_M4 0.035
r 32000_60000_M3 32000_60000_M4 0.035
r 32000_64000_M3 32000_64000_M4 0.035
r 32000_68000_M3 32000_68000_M4 0.035
r 32000_72000_M3 32000_72000_M4 0.035
r 32000_76000_M3 32000_76000_M4 0.035
r 32000_80000_M3 32000_80000_M4 0.035
r 32000_84000_M3 32000_84000_M4 0.035
r 32000_88000_M3 32000_88000_M4 0.035
r 32000_92000_M3 32000_92000_M4 0.035
r 32000_96000_M3 32000_96000_M4 0.035
r 32000_100000_M3 32000_100000_M4 0.035
r 36000_4000_M3 36000_4000_M4 0.035
r 36000_8000_M3 36000_8000_M4 0.035
r 36000_12000_M3 36000_12000_M4 0.035
r 36000_16000_M3 36000_16000_M4 0.035
r 36000_20000_M3 36000_20000_M4 0.035
r 36000_24000_M3 36000_24000_M4 0.035
r 36000_28000_M3 36000_28000_M4 0.035
r 36000_32000_M3 36000_32000_M4 0.035
r 36000_36000_M3 36000_36000_M4 0.035
r 36000_40000_M3 36000_40000_M4 0.035
r 36000_44000_M3 36000_44000_M4 0.035
r 36000_48000_M3 36000_48000_M4 0.035
r 36000_52000_M3 36000_52000_M4 0.035
r 36000_56000_M3 36000_56000_M4 0.035
r 36000_60000_M3 36000_60000_M4 0.035
r 36000_64000_M3 36000_64000_M4 0.035
r 36000_68000_M3 36000_68000_M4 0.035
r 36000_72000_M3 36000_72000_M4 0.035
r 36000_76000_M3 36000_76000_M4 0.035
r 36000_80000_M3 36000_80000_M4 0.035
r 36000_84000_M3 36000_84000_M4 0.035
r 36000_88000_M3 36000_88000_M4 0.035
r 36000_92000_M3 36000_92000_M4 0.035
r 36000_96000_M3 36000_96000_M4 0.035
r 36000_100000_M3 36000_100000_M4 0.035
r 40000_4000_M3 40000_4000_M4 0.035
r 40000_8000_M3 40000_8000_M4 0.035
r 40000_12000_M3 40000_12000_M4 0.035
r 40000_16000_M3 40000_16000_M4 0.035
r 40000_20000_M3 40000_20000_M4 0.035
r 40000_24000_M3 40000_24000_M4 0.035
r 40000_28000_M3 40000_28000_M4 0.035
r 40000_32000_M3 40000_32000_M4 0.035
r 40000_36000_M3 40000_36000_M4 0.035
r 40000_40000_M3 40000_40000_M4 0.035
r 40000_44000_M3 40000_44000_M4 0.035
r 40000_48000_M3 40000_48000_M4 0.035
r 40000_52000_M3 40000_52000_M4 0.035
r 40000_56000_M3 40000_56000_M4 0.035
r 40000_60000_M3 40000_60000_M4 0.035
r 40000_64000_M3 40000_64000_M4 0.035
r 40000_68000_M3 40000_68000_M4 0.035
r 40000_72000_M3 40000_72000_M4 0.035
r 40000_76000_M3 40000_76000_M4 0.035
r 40000_80000_M3 40000_80000_M4 0.035
r 40000_84000_M3 40000_84000_M4 0.035
r 40000_88000_M3 40000_88000_M4 0.035
r 40000_92000_M3 40000_92000_M4 0.035
r 40000_96000_M3 40000_96000_M4 0.035
r 40000_100000_M3 40000_100000_M4 0.035
r 44000_4000_M3 44000_4000_M4 0.035
r 44000_8000_M3 44000_8000_M4 0.035
r 44000_12000_M3 44000_12000_M4 0.035
r 44000_16000_M3 44000_16000_M4 0.035
r 44000_20000_M3 44000_20000_M4 0.035
r 44000_24000_M3 44000_24000_M4 0.035
r 44000_28000_M3 44000_28000_M4 0.035
r 44000_32000_M3 44000_32000_M4 0.035
r 44000_36000_M3 44000_36000_M4 0.035
r 44000_40000_M3 44000_40000_M4 0.035
r 44000_44000_M3 44000_44000_M4 0.035
r 44000_48000_M3 44000_48000_M4 0.035
r 44000_52000_M3 44000_52000_M4 0.035
r 44000_56000_M3 44000_56000_M4 0.035
r 44000_60000_M3 44000_60000_M4 0.035
r 44000_64000_M3 44000_64000_M4 0.035
r 44000_68000_M3 44000_68000_M4 0.035
r 44000_72000_M3 44000_72000_M4 0.035
r 44000_76000_M3 44000_76000_M4 0.035
r 44000_80000_M3 44000_80000_M4 0.035
r 44000_84000_M3 44000_84000_M4 0.035
r 44000_88000_M3 44000_88000_M4 0.035
r 44000_92000_M3 44000_92000_M4 0.035
r 44000_96000_M3 44000_96000_M4 0.035
r 44000_100000_M3 44000_100000_M4 0.035
r 48000_4000_M3 48000_4000_M4 0.035
r 48000_8000_M3 48000_8000_M4 0.035
r 48000_12000_M3 48000_12000_M4 0.035
r 48000_16000_M3 48000_16000_M4 0.035
r 48000_20000_M3 48000_20000_M4 0.035
r 48000_24000_M3 48000_24000_M4 0.035
r 48000_28000_M3 48000_28000_M4 0.035
r 48000_32000_M3 48000_32000_M4 0.035
r 48000_36000_M3 48000_36000_M4 0.035
r 48000_40000_M3 48000_40000_M4 0.035
r 48000_44000_M3 48000_44000_M4 0.035
r 48000_48000_M3 48000_48000_M4 0.035
r 48000_52000_M3 48000_52000_M4 0.035
r 48000_56000_M3 48000_56000_M4 0.035
r 48000_60000_M3 48000_60000_M4 0.035
r 48000_64000_M3 48000_64000_M4 0.035
r 48000_68000_M3 48000_68000_M4 0.035
r 48000_72000_M3 48000_72000_M4 0.035
r 48000_76000_M3 48000_76000_M4 0.035
r 48000_80000_M3 48000_80000_M4 0.035
r 48000_84000_M3 48000_84000_M4 0.035
r 48000_88000_M3 48000_88000_M4 0.035
r 48000_92000_M3 48000_92000_M4 0.035
r 48000_96000_M3 48000_96000_M4 0.035
r 48000_100000_M3 48000_100000_M4 0.035
r 52000_4000_M3 52000_4000_M4 0.035
r 52000_8000_M3 52000_8000_M4 0.035
r 52000_12000_M3 52000_12000_M4 0.035
r 52000_16000_M3 52000_16000_M4 0.035
r 52000_20000_M3 52000_20000_M4 0.035
r 52000_24000_M3 52000_24000_M4 0.035
r 52000_28000_M3 52000_28000_M4 0.035
r 52000_32000_M3 52000_32000_M4 0.035
r 52000_36000_M3 52000_36000_M4 0.035
r 52000_40000_M3 52000_40000_M4 0.035
r 52000_44000_M3 52000_44000_M4 0.035
r 52000_48000_M3 52000_48000_M4 0.035
r 52000_52000_M3 52000_52000_M4 0.035
r 52000_56000_M3 52000_56000_M4 0.035
r 52000_60000_M3 52000_60000_M4 0.035
r 52000_64000_M3 52000_64000_M4 0.035
r 52000_68000_M3 52000_68000_M4 0.035
r 52000_72000_M3 52000_72000_M4 0.035
r 52000_76000_M3 52000_76000_M4 0.035
r 52000_80000_M3 52000_80000_M4 0.035
r 52000_84000_M3 52000_84000_M4 0.035
r 52000_88000_M3 52000_88000_M4 0.035
r 52000_92000_M3 52000_92000_M4 0.035
r 52000_96000_M3 52000_96000_M4 0.035
r 52000_100000_M3 52000_100000_M4 0.035
r 56000_4000_M3 56000_4000_M4 0.035
r 56000_8000_M3 56000_8000_M4 0.035
r 56000_12000_M3 56000_12000_M4 0.035
r 56000_16000_M3 56000_16000_M4 0.035
r 56000_20000_M3 56000_20000_M4 0.035
r 56000_24000_M3 56000_24000_M4 0.035
r 56000_28000_M3 56000_28000_M4 0.035
r 56000_32000_M3 56000_32000_M4 0.035
r 56000_36000_M3 56000_36000_M4 0.035
r 56000_40000_M3 56000_40000_M4 0.035
r 56000_44000_M3 56000_44000_M4 0.035
r 56000_48000_M3 56000_48000_M4 0.035
r 56000_52000_M3 56000_52000_M4 0.035
r 56000_56000_M3 56000_56000_M4 0.035
r 56000_60000_M3 56000_60000_M4 0.035
r 56000_64000_M3 56000_64000_M4 0.035
r 56000_68000_M3 56000_68000_M4 0.035
r 56000_72000_M3 56000_72000_M4 0.035
r 56000_76000_M3 56000_76000_M4 0.035
r 56000_80000_M3 56000_80000_M4 0.035
r 56000_84000_M3 56000_84000_M4 0.035
r 56000_88000_M3 56000_88000_M4 0.035
r 56000_92000_M3 56000_92000_M4 0.035
r 56000_96000_M3 56000_96000_M4 0.035
r 56000_100000_M3 56000_100000_M4 0.035
r 60000_4000_M3 60000_4000_M4 0.035
r 60000_8000_M3 60000_8000_M4 0.035
r 60000_12000_M3 60000_12000_M4 0.035
r 60000_16000_M3 60000_16000_M4 0.035
r 60000_20000_M3 60000_20000_M4 0.035
r 60000_24000_M3 60000_24000_M4 0.035
r 60000_28000_M3 60000_28000_M4 0.035
r 60000_32000_M3 60000_32000_M4 0.035
r 60000_36000_M3 60000_36000_M4 0.035
r 60000_40000_M3 60000_40000_M4 0.035
r 60000_44000_M3 60000_44000_M4 0.035
r 60000_48000_M3 60000_48000_M4 0.035
r 60000_52000_M3 60000_52000_M4 0.035
r 60000_56000_M3 60000_56000_M4 0.035
r 60000_60000_M3 60000_60000_M4 0.035
r 60000_64000_M3 60000_64000_M4 0.035
r 60000_68000_M3 60000_68000_M4 0.035
r 60000_72000_M3 60000_72000_M4 0.035
r 60000_76000_M3 60000_76000_M4 0.035
r 60000_80000_M3 60000_80000_M4 0.035
r 60000_84000_M3 60000_84000_M4 0.035
r 60000_88000_M3 60000_88000_M4 0.035
r 60000_92000_M3 60000_92000_M4 0.035
r 60000_96000_M3 60000_96000_M4 0.035
r 60000_100000_M3 60000_100000_M4 0.035
r 64000_4000_M3 64000_4000_M4 0.035
r 64000_8000_M3 64000_8000_M4 0.035
r 64000_12000_M3 64000_12000_M4 0.035
r 64000_16000_M3 64000_16000_M4 0.035
r 64000_20000_M3 64000_20000_M4 0.035
r 64000_24000_M3 64000_24000_M4 0.035
r 64000_28000_M3 64000_28000_M4 0.035
r 64000_32000_M3 64000_32000_M4 0.035
r 64000_36000_M3 64000_36000_M4 0.035
r 64000_40000_M3 64000_40000_M4 0.035
r 64000_44000_M3 64000_44000_M4 0.035
r 64000_48000_M3 64000_48000_M4 0.035
r 64000_52000_M3 64000_52000_M4 0.035
r 64000_56000_M3 64000_56000_M4 0.035
r 64000_60000_M3 64000_60000_M4 0.035
r 64000_64000_M3 64000_64000_M4 0.035
r 64000_68000_M3 64000_68000_M4 0.035
r 64000_72000_M3 64000_72000_M4 0.035
r 64000_76000_M3 64000_76000_M4 0.035
r 64000_80000_M3 64000_80000_M4 0.035
r 64000_84000_M3 64000_84000_M4 0.035
r 64000_88000_M3 64000_88000_M4 0.035
r 64000_92000_M3 64000_92000_M4 0.035
r 64000_96000_M3 64000_96000_M4 0.035
r 64000_100000_M3 64000_100000_M4 0.035
r 68000_4000_M3 68000_4000_M4 0.035
r 68000_8000_M3 68000_8000_M4 0.035
r 68000_12000_M3 68000_12000_M4 0.035
r 68000_16000_M3 68000_16000_M4 0.035
r 68000_20000_M3 68000_20000_M4 0.035
r 68000_24000_M3 68000_24000_M4 0.035
r 68000_28000_M3 68000_28000_M4 0.035
r 68000_32000_M3 68000_32000_M4 0.035
r 68000_36000_M3 68000_36000_M4 0.035
r 68000_40000_M3 68000_40000_M4 0.035
r 68000_44000_M3 68000_44000_M4 0.035
r 68000_48000_M3 68000_48000_M4 0.035
r 68000_52000_M3 68000_52000_M4 0.035
r 68000_56000_M3 68000_56000_M4 0.035
r 68000_60000_M3 68000_60000_M4 0.035
r 68000_64000_M3 68000_64000_M4 0.035
r 68000_68000_M3 68000_68000_M4 0.035
r 68000_72000_M3 68000_72000_M4 0.035
r 68000_76000_M3 68000_76000_M4 0.035
r 68000_80000_M3 68000_80000_M4 0.035
r 68000_84000_M3 68000_84000_M4 0.035
r 68000_88000_M3 68000_88000_M4 0.035
r 68000_92000_M3 68000_92000_M4 0.035
r 68000_96000_M3 68000_96000_M4 0.035
r 68000_100000_M3 68000_100000_M4 0.035
r 72000_4000_M3 72000_4000_M4 0.035
r 72000_8000_M3 72000_8000_M4 0.035
r 72000_12000_M3 72000_12000_M4 0.035
r 72000_16000_M3 72000_16000_M4 0.035
r 72000_20000_M3 72000_20000_M4 0.035
r 72000_24000_M3 72000_24000_M4 0.035
r 72000_28000_M3 72000_28000_M4 0.035
r 72000_32000_M3 72000_32000_M4 0.035
r 72000_36000_M3 72000_36000_M4 0.035
r 72000_40000_M3 72000_40000_M4 0.035
r 72000_44000_M3 72000_44000_M4 0.035
r 72000_48000_M3 72000_48000_M4 0.035
r 72000_52000_M3 72000_52000_M4 0.035
r 72000_56000_M3 72000_56000_M4 0.035
r 72000_60000_M3 72000_60000_M4 0.035
r 72000_64000_M3 72000_64000_M4 0.035
r 72000_68000_M3 72000_68000_M4 0.035
r 72000_72000_M3 72000_72000_M4 0.035
r 72000_76000_M3 72000_76000_M4 0.035
r 72000_80000_M3 72000_80000_M4 0.035
r 72000_84000_M3 72000_84000_M4 0.035
r 72000_88000_M3 72000_88000_M4 0.035
r 72000_92000_M3 72000_92000_M4 0.035
r 72000_96000_M3 72000_96000_M4 0.035
r 72000_100000_M3 72000_100000_M4 0.035
r 76000_4000_M3 76000_4000_M4 0.035
r 76000_8000_M3 76000_8000_M4 0.035
r 76000_12000_M3 76000_12000_M4 0.035
r 76000_16000_M3 76000_16000_M4 0.035
r 76000_20000_M3 76000_20000_M4 0.035
r 76000_24000_M3 76000_24000_M4 0.035
r 76000_28000_M3 76000_28000_M4 0.035
r 76000_32000_M3 76000_32000_M4 0.035
r 76000_36000_M3 76000_36000_M4 0.035
r 76000_40000_M3 76000_40000_M4 0.035
r 76000_44000_M3 76000_44000_M4 0.035
r 76000_48000_M3 76000_48000_M4 0.035
r 76000_52000_M3 76000_52000_M4 0.035
r 76000_56000_M3 76000_56000_M4 0.035
r 76000_60000_M3 76000_60000_M4 0.035
r 76000_64000_M3 76000_64000_M4 0.035
r 76000_68000_M3 76000_68000_M4 0.035
r 76000_72000_M3 76000_72000_M4 0.035
r 76000_76000_M3 76000_76000_M4 0.035
r 76000_80000_M3 76000_80000_M4 0.035
r 76000_84000_M3 76000_84000_M4 0.035
r 76000_88000_M3 76000_88000_M4 0.035
r 76000_92000_M3 76000_92000_M4 0.035
r 76000_96000_M3 76000_96000_M4 0.035
r 76000_100000_M3 76000_100000_M4 0.035
r 80000_4000_M3 80000_4000_M4 0.035
r 80000_8000_M3 80000_8000_M4 0.035
r 80000_12000_M3 80000_12000_M4 0.035
r 80000_16000_M3 80000_16000_M4 0.035
r 80000_20000_M3 80000_20000_M4 0.035
r 80000_24000_M3 80000_24000_M4 0.035
r 80000_28000_M3 80000_28000_M4 0.035
r 80000_32000_M3 80000_32000_M4 0.035
r 80000_36000_M3 80000_36000_M4 0.035
r 80000_40000_M3 80000_40000_M4 0.035
r 80000_44000_M3 80000_44000_M4 0.035
r 80000_48000_M3 80000_48000_M4 0.035
r 80000_52000_M3 80000_52000_M4 0.035
r 80000_56000_M3 80000_56000_M4 0.035
r 80000_60000_M3 80000_60000_M4 0.035
r 80000_64000_M3 80000_64000_M4 0.035
r 80000_68000_M3 80000_68000_M4 0.035
r 80000_72000_M3 80000_72000_M4 0.035
r 80000_76000_M3 80000_76000_M4 0.035
r 80000_80000_M3 80000_80000_M4 0.035
r 80000_84000_M3 80000_84000_M4 0.035
r 80000_88000_M3 80000_88000_M4 0.035
r 80000_92000_M3 80000_92000_M4 0.035
r 80000_96000_M3 80000_96000_M4 0.035
r 80000_100000_M3 80000_100000_M4 0.035
r 84000_4000_M3 84000_4000_M4 0.035
r 84000_8000_M3 84000_8000_M4 0.035
r 84000_12000_M3 84000_12000_M4 0.035
r 84000_16000_M3 84000_16000_M4 0.035
r 84000_20000_M3 84000_20000_M4 0.035
r 84000_24000_M3 84000_24000_M4 0.035
r 84000_28000_M3 84000_28000_M4 0.035
r 84000_32000_M3 84000_32000_M4 0.035
r 84000_36000_M3 84000_36000_M4 0.035
r 84000_40000_M3 84000_40000_M4 0.035
r 84000_44000_M3 84000_44000_M4 0.035
r 84000_48000_M3 84000_48000_M4 0.035
r 84000_52000_M3 84000_52000_M4 0.035
r 84000_56000_M3 84000_56000_M4 0.035
r 84000_60000_M3 84000_60000_M4 0.035
r 84000_64000_M3 84000_64000_M4 0.035
r 84000_68000_M3 84000_68000_M4 0.035
r 84000_72000_M3 84000_72000_M4 0.035
r 84000_76000_M3 84000_76000_M4 0.035
r 84000_80000_M3 84000_80000_M4 0.035
r 84000_84000_M3 84000_84000_M4 0.035
r 84000_88000_M3 84000_88000_M4 0.035
r 84000_92000_M3 84000_92000_M4 0.035
r 84000_96000_M3 84000_96000_M4 0.035
r 84000_100000_M3 84000_100000_M4 0.035
r 88000_4000_M3 88000_4000_M4 0.035
r 88000_8000_M3 88000_8000_M4 0.035
r 88000_12000_M3 88000_12000_M4 0.035
r 88000_16000_M3 88000_16000_M4 0.035
r 88000_20000_M3 88000_20000_M4 0.035
r 88000_24000_M3 88000_24000_M4 0.035
r 88000_28000_M3 88000_28000_M4 0.035
r 88000_32000_M3 88000_32000_M4 0.035
r 88000_36000_M3 88000_36000_M4 0.035
r 88000_40000_M3 88000_40000_M4 0.035
r 88000_44000_M3 88000_44000_M4 0.035
r 88000_48000_M3 88000_48000_M4 0.035
r 88000_52000_M3 88000_52000_M4 0.035
r 88000_56000_M3 88000_56000_M4 0.035
r 88000_60000_M3 88000_60000_M4 0.035
r 88000_64000_M3 88000_64000_M4 0.035
r 88000_68000_M3 88000_68000_M4 0.035
r 88000_72000_M3 88000_72000_M4 0.035
r 88000_76000_M3 88000_76000_M4 0.035
r 88000_80000_M3 88000_80000_M4 0.035
r 88000_84000_M3 88000_84000_M4 0.035
r 88000_88000_M3 88000_88000_M4 0.035
r 88000_92000_M3 88000_92000_M4 0.035
r 88000_96000_M3 88000_96000_M4 0.035
r 88000_100000_M3 88000_100000_M4 0.035
r 92000_4000_M3 92000_4000_M4 0.035
r 92000_8000_M3 92000_8000_M4 0.035
r 92000_12000_M3 92000_12000_M4 0.035
r 92000_16000_M3 92000_16000_M4 0.035
r 92000_20000_M3 92000_20000_M4 0.035
r 92000_24000_M3 92000_24000_M4 0.035
r 92000_28000_M3 92000_28000_M4 0.035
r 92000_32000_M3 92000_32000_M4 0.035
r 92000_36000_M3 92000_36000_M4 0.035
r 92000_40000_M3 92000_40000_M4 0.035
r 92000_44000_M3 92000_44000_M4 0.035
r 92000_48000_M3 92000_48000_M4 0.035
r 92000_52000_M3 92000_52000_M4 0.035
r 92000_56000_M3 92000_56000_M4 0.035
r 92000_60000_M3 92000_60000_M4 0.035
r 92000_64000_M3 92000_64000_M4 0.035
r 92000_68000_M3 92000_68000_M4 0.035
r 92000_72000_M3 92000_72000_M4 0.035
r 92000_76000_M3 92000_76000_M4 0.035
r 92000_80000_M3 92000_80000_M4 0.035
r 92000_84000_M3 92000_84000_M4 0.035
r 92000_88000_M3 92000_88000_M4 0.035
r 92000_92000_M3 92000_92000_M4 0.035
r 92000_96000_M3 92000_96000_M4 0.035
r 92000_100000_M3 92000_100000_M4 0.035
r 96000_4000_M3 96000_4000_M4 0.035
r 96000_8000_M3 96000_8000_M4 0.035
r 96000_12000_M3 96000_12000_M4 0.035
r 96000_16000_M3 96000_16000_M4 0.035
r 96000_20000_M3 96000_20000_M4 0.035
r 96000_24000_M3 96000_24000_M4 0.035
r 96000_28000_M3 96000_28000_M4 0.035
r 96000_32000_M3 96000_32000_M4 0.035
r 96000_36000_M3 96000_36000_M4 0.035
r 96000_40000_M3 96000_40000_M4 0.035
r 96000_44000_M3 96000_44000_M4 0.035
r 96000_48000_M3 96000_48000_M4 0.035
r 96000_52000_M3 96000_52000_M4 0.035
r 96000_56000_M3 96000_56000_M4 0.035
r 96000_60000_M3 96000_60000_M4 0.035
r 96000_64000_M3 96000_64000_M4 0.035
r 96000_68000_M3 96000_68000_M4 0.035
r 96000_72000_M3 96000_72000_M4 0.035
r 96000_76000_M3 96000_76000_M4 0.035
r 96000_80000_M3 96000_80000_M4 0.035
r 96000_84000_M3 96000_84000_M4 0.035
r 96000_88000_M3 96000_88000_M4 0.035
r 96000_92000_M3 96000_92000_M4 0.035
r 96000_96000_M3 96000_96000_M4 0.035
r 96000_100000_M3 96000_100000_M4 0.035
r 100000_4000_M3 100000_4000_M4 0.035
r 100000_8000_M3 100000_8000_M4 0.035
r 100000_12000_M3 100000_12000_M4 0.035
r 100000_16000_M3 100000_16000_M4 0.035
r 100000_20000_M3 100000_20000_M4 0.035
r 100000_24000_M3 100000_24000_M4 0.035
r 100000_28000_M3 100000_28000_M4 0.035
r 100000_32000_M3 100000_32000_M4 0.035
r 100000_36000_M3 100000_36000_M4 0.035
r 100000_40000_M3 100000_40000_M4 0.035
r 100000_44000_M3 100000_44000_M4 0.035
r 100000_48000_M3 100000_48000_M4 0.035
r 100000_52000_M3 100000_52000_M4 0.035
r 100000_56000_M3 100000_56000_M4 0.035
r 100000_60000_M3 100000_60000_M4 0.035
r 100000_64000_M3 100000_64000_M4 0.035
r 100000_68000_M3 100000_68000_M4 0.035
r 100000_72000_M3 100000_72000_M4 0.035
r 100000_76000_M3 100000_76000_M4 0.035
r 100000_80000_M3 100000_80000_M4 0.035
r 100000_84000_M3 100000_84000_M4 0.035
r 100000_88000_M3 100000_88000_M4 0.035
r 100000_92000_M3 100000_92000_M4 0.035
r 100000_96000_M3 100000_96000_M4 0.035
r 100000_100000_M3 100000_100000_M4 0.035

* ============================================================================
* Via connections M4 to M5
* ============================================================================

r 8000_8000_M4 8000_8000_M5 0.030
r 8000_16000_M4 8000_16000_M5 0.030
r 8000_24000_M4 8000_24000_M5 0.030
r 8000_32000_M4 8000_32000_M5 0.030
r 8000_40000_M4 8000_40000_M5 0.030
r 8000_48000_M4 8000_48000_M5 0.030
r 8000_56000_M4 8000_56000_M5 0.030
r 8000_64000_M4 8000_64000_M5 0.030
r 8000_72000_M4 8000_72000_M5 0.030
r 8000_80000_M4 8000_80000_M5 0.030
r 8000_88000_M4 8000_88000_M5 0.030
r 8000_96000_M4 8000_96000_M5 0.030
r 16000_8000_M4 16000_8000_M5 0.030
r 16000_16000_M4 16000_16000_M5 0.030
r 16000_24000_M4 16000_24000_M5 0.030
r 16000_32000_M4 16000_32000_M5 0.030
r 16000_40000_M4 16000_40000_M5 0.030
r 16000_48000_M4 16000_48000_M5 0.030
r 16000_56000_M4 16000_56000_M5 0.030
r 16000_64000_M4 16000_64000_M5 0.030
r 16000_72000_M4 16000_72000_M5 0.030
r 16000_80000_M4 16000_80000_M5 0.030
r 16000_88000_M4 16000_88000_M5 0.030
r 16000_96000_M4 16000_96000_M5 0.030
r 24000_8000_M4 24000_8000_M5 0.030
r 24000_16000_M4 24000_16000_M5 0.030
r 24000_24000_M4 24000_24000_M5 0.030
r 24000_32000_M4 24000_32000_M5 0.030
r 24000_40000_M4 24000_40000_M5 0.030
r 24000_48000_M4 24000_48000_M5 0.030
r 24000_56000_M4 24000_56000_M5 0.030
r 24000_64000_M4 24000_64000_M5 0.030
r 24000_72000_M4 24000_72000_M5 0.030
r 24000_80000_M4 24000_80000_M5 0.030
r 24000_88000_M4 24000_88000_M5 0.030
r 24000_96000_M4 24000_96000_M5 0.030
r 32000_8000_M4 32000_8000_M5 0.030
r 32000_16000_M4 32000_16000_M5 0.030
r 32000_24000_M4 32000_24000_M5 0.030
r 32000_32000_M4 32000_32000_M5 0.030
r 32000_40000_M4 32000_40000_M5 0.030
r 32000_48000_M4 32000_48000_M5 0.030
r 32000_56000_M4 32000_56000_M5 0.030
r 32000_64000_M4 32000_64000_M5 0.030
r 32000_72000_M4 32000_72000_M5 0.030
r 32000_80000_M4 32000_80000_M5 0.030
r 32000_88000_M4 32000_88000_M5 0.030
r 32000_96000_M4 32000_96000_M5 0.030
r 40000_8000_M4 40000_8000_M5 0.030
r 40000_16000_M4 40000_16000_M5 0.030
r 40000_24000_M4 40000_24000_M5 0.030
r 40000_32000_M4 40000_32000_M5 0.030
r 40000_40000_M4 40000_40000_M5 0.030
r 40000_48000_M4 40000_48000_M5 0.030
r 40000_56000_M4 40000_56000_M5 0.030
r 40000_64000_M4 40000_64000_M5 0.030
r 40000_72000_M4 40000_72000_M5 0.030
r 40000_80000_M4 40000_80000_M5 0.030
r 40000_88000_M4 40000_88000_M5 0.030
r 40000_96000_M4 40000_96000_M5 0.030
r 48000_8000_M4 48000_8000_M5 0.030
r 48000_16000_M4 48000_16000_M5 0.030
r 48000_24000_M4 48000_24000_M5 0.030
r 48000_32000_M4 48000_32000_M5 0.030
r 48000_40000_M4 48000_40000_M5 0.030
r 48000_48000_M4 48000_48000_M5 0.030
r 48000_56000_M4 48000_56000_M5 0.030
r 48000_64000_M4 48000_64000_M5 0.030
r 48000_72000_M4 48000_72000_M5 0.030
r 48000_80000_M4 48000_80000_M5 0.030
r 48000_88000_M4 48000_88000_M5 0.030
r 48000_96000_M4 48000_96000_M5 0.030
r 56000_8000_M4 56000_8000_M5 0.030
r 56000_16000_M4 56000_16000_M5 0.030
r 56000_24000_M4 56000_24000_M5 0.030
r 56000_32000_M4 56000_32000_M5 0.030
r 56000_40000_M4 56000_40000_M5 0.030
r 56000_48000_M4 56000_48000_M5 0.030
r 56000_56000_M4 56000_56000_M5 0.030
r 56000_64000_M4 56000_64000_M5 0.030
r 56000_72000_M4 56000_72000_M5 0.030
r 56000_80000_M4 56000_80000_M5 0.030
r 56000_88000_M4 56000_88000_M5 0.030
r 56000_96000_M4 56000_96000_M5 0.030
r 64000_8000_M4 64000_8000_M5 0.030
r 64000_16000_M4 64000_16000_M5 0.030
r 64000_24000_M4 64000_24000_M5 0.030
r 64000_32000_M4 64000_32000_M5 0.030
r 64000_40000_M4 64000_40000_M5 0.030
r 64000_48000_M4 64000_48000_M5 0.030
r 64000_56000_M4 64000_56000_M5 0.030
r 64000_64000_M4 64000_64000_M5 0.030
r 64000_72000_M4 64000_72000_M5 0.030
r 64000_80000_M4 64000_80000_M5 0.030
r 64000_88000_M4 64000_88000_M5 0.030
r 64000_96000_M4 64000_96000_M5 0.030
r 72000_8000_M4 72000_8000_M5 0.030
r 72000_16000_M4 72000_16000_M5 0.030
r 72000_24000_M4 72000_24000_M5 0.030
r 72000_32000_M4 72000_32000_M5 0.030
r 72000_40000_M4 72000_40000_M5 0.030
r 72000_48000_M4 72000_48000_M5 0.030
r 72000_56000_M4 72000_56000_M5 0.030
r 72000_64000_M4 72000_64000_M5 0.030
r 72000_72000_M4 72000_72000_M5 0.030
r 72000_80000_M4 72000_80000_M5 0.030
r 72000_88000_M4 72000_88000_M5 0.030
r 72000_96000_M4 72000_96000_M5 0.030
r 80000_8000_M4 80000_8000_M5 0.030
r 80000_16000_M4 80000_16000_M5 0.030
r 80000_24000_M4 80000_24000_M5 0.030
r 80000_32000_M4 80000_32000_M5 0.030
r 80000_40000_M4 80000_40000_M5 0.030
r 80000_48000_M4 80000_48000_M5 0.030
r 80000_56000_M4 80000_56000_M5 0.030
r 80000_64000_M4 80000_64000_M5 0.030
r 80000_72000_M4 80000_72000_M5 0.030
r 80000_80000_M4 80000_80000_M5 0.030
r 80000_88000_M4 80000_88000_M5 0.030
r 80000_96000_M4 80000_96000_M5 0.030
r 88000_8000_M4 88000_8000_M5 0.030
r 88000_16000_M4 88000_16000_M5 0.030
r 88000_24000_M4 88000_24000_M5 0.030
r 88000_32000_M4 88000_32000_M5 0.030
r 88000_40000_M4 88000_40000_M5 0.030
r 88000_48000_M4 88000_48000_M5 0.030
r 88000_56000_M4 88000_56000_M5 0.030
r 88000_64000_M4 88000_64000_M5 0.030
r 88000_72000_M4 88000_72000_M5 0.030
r 88000_80000_M4 88000_80000_M5 0.030
r 88000_88000_M4 88000_88000_M5 0.030
r 88000_96000_M4 88000_96000_M5 0.030
r 96000_8000_M4 96000_8000_M5 0.030
r 96000_16000_M4 96000_16000_M5 0.030
r 96000_24000_M4 96000_24000_M5 0.030
r 96000_32000_M4 96000_32000_M5 0.030
r 96000_40000_M4 96000_40000_M5 0.030
r 96000_48000_M4 96000_48000_M5 0.030
r 96000_56000_M4 96000_56000_M5 0.030
r 96000_64000_M4 96000_64000_M5 0.030
r 96000_72000_M4 96000_72000_M5 0.030
r 96000_80000_M4 96000_80000_M5 0.030
r 96000_88000_M4 96000_88000_M5 0.030
r 96000_96000_M4 96000_96000_M5 0.030

* ============================================================================
* ISOLATED ISLANDS - Not connected to main grid
* These test floating/disconnected load handling
* ============================================================================

* island1: 3x3 grid at (110000, 10000)
r 110000_10000_M1 112000_10000_M1 0.020
r 112000_10000_M1 114000_10000_M1 0.020
r 110000_12000_M1 112000_12000_M1 0.020
r 112000_12000_M1 114000_12000_M1 0.020
r 110000_14000_M1 112000_14000_M1 0.020
r 112000_14000_M1 114000_14000_M1 0.020
r 110000_10000_M1 110000_12000_M1 0.025
r 110000_12000_M1 110000_14000_M1 0.025
r 112000_10000_M1 112000_12000_M1 0.025
r 112000_12000_M1 112000_14000_M1 0.025
r 114000_10000_M1 114000_12000_M1 0.025
r 114000_12000_M1 114000_14000_M1 0.025

* island2: 3x3 grid at (110000, 30000)
r 110000_30000_M1 112000_30000_M1 0.020
r 112000_30000_M1 114000_30000_M1 0.020
r 110000_32000_M1 112000_32000_M1 0.020
r 112000_32000_M1 114000_32000_M1 0.020
r 110000_34000_M1 112000_34000_M1 0.020
r 112000_34000_M1 114000_34000_M1 0.020
r 110000_30000_M1 110000_32000_M1 0.025
r 110000_32000_M1 110000_34000_M1 0.025
r 112000_30000_M1 112000_32000_M1 0.025
r 112000_32000_M1 112000_34000_M1 0.025
r 114000_30000_M1 114000_32000_M1 0.025
r 114000_32000_M1 114000_34000_M1 0.025

* island3: 4x4 grid at (110000, 50000)
r 110000_50000_M1 112000_50000_M1 0.020
r 112000_50000_M1 114000_50000_M1 0.020
r 114000_50000_M1 116000_50000_M1 0.020
r 110000_52000_M1 112000_52000_M1 0.020
r 112000_52000_M1 114000_52000_M1 0.020
r 114000_52000_M1 116000_52000_M1 0.020
r 110000_54000_M1 112000_54000_M1 0.020
r 112000_54000_M1 114000_54000_M1 0.020
r 114000_54000_M1 116000_54000_M1 0.020
r 110000_56000_M1 112000_56000_M1 0.020
r 112000_56000_M1 114000_56000_M1 0.020
r 114000_56000_M1 116000_56000_M1 0.020
r 110000_50000_M1 110000_52000_M1 0.025
r 110000_52000_M1 110000_54000_M1 0.025
r 110000_54000_M1 110000_56000_M1 0.025
r 112000_50000_M1 112000_52000_M1 0.025
r 112000_52000_M1 112000_54000_M1 0.025
r 112000_54000_M1 112000_56000_M1 0.025
r 114000_50000_M1 114000_52000_M1 0.025
r 114000_52000_M1 114000_54000_M1 0.025
r 114000_54000_M1 114000_56000_M1 0.025
r 116000_50000_M1 116000_52000_M1 0.025
r 116000_52000_M1 116000_54000_M1 0.025
r 116000_54000_M1 116000_56000_M1 0.025