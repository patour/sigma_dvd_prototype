* Tile 0_0 - Die resistor/capacitor mesh
* Two-layer structure: M1 (horizontal stripes) and M2 (vertical stripes)
* 5x5 grid on each layer with via connections

* ============================================================================
* Layer M1 - Horizontal routing (5 rows)
* ============================================================================

* Row 1 (y=1000)
r 1000_1000_M1 2000_1000_M1 0.020
r 2000_1000_M1 3000_1000_M1 0.020
r 3000_1000_M1 4000_1000_M1 0.020
r 4000_1000_M1 5000_1000_M1 0.020

* Row 2 (y=2000)
r 1000_2000_M1 2000_2000_M1 0.020
r 2000_2000_M1 3000_2000_M1 0.020
r 3000_2000_M1 4000_2000_M1 0.020
r 4000_2000_M1 5000_2000_M1 0.020

* Row 3 (y=3000)
r 1000_3000_M1 2000_3000_M1 0.020
r 2000_3000_M1 3000_3000_M1 0.020
r 3000_3000_M1 4000_3000_M1 0.020
r 4000_3000_M1 5000_3000_M1 0.020

* Row 4 (y=4000)
r 1000_4000_M1 2000_4000_M1 0.020
r 2000_4000_M1 3000_4000_M1 0.020
r 3000_4000_M1 4000_4000_M1 0.020
r 4000_4000_M1 5000_4000_M1 0.020

* Row 5 (y=5000)
r 1000_5000_M1 2000_5000_M1 0.020
r 2000_5000_M1 3000_5000_M1 0.020
r 3000_5000_M1 4000_5000_M1 0.020
r 4000_5000_M1 5000_5000_M1 0.020

* ============================================================================
* Layer M2 - Vertical routing (5 columns)
* ============================================================================

* Column 1 (x=1000)
r 1000_1000_M2 1000_2000_M2 0.015
r 1000_2000_M2 1000_3000_M2 0.015
r 1000_3000_M2 1000_4000_M2 0.015
r 1000_4000_M2 1000_5000_M2 0.015

* Column 2 (x=2000)
r 2000_1000_M2 2000_2000_M2 0.015
r 2000_2000_M2 2000_3000_M2 0.015
r 2000_3000_M2 2000_4000_M2 0.015
r 2000_4000_M2 2000_5000_M2 0.015

* Column 3 (x=3000)
r 3000_1000_M2 3000_2000_M2 0.015
r 3000_2000_M2 3000_3000_M2 0.015
r 3000_3000_M2 3000_4000_M2 0.015
r 3000_4000_M2 3000_5000_M2 0.015

* Column 4 (x=4000)
r 4000_1000_M2 4000_2000_M2 0.015
r 4000_2000_M2 4000_3000_M2 0.015
r 4000_3000_M2 4000_4000_M2 0.015
r 4000_4000_M2 4000_5000_M2 0.015

* Column 5 (x=5000)
r 5000_1000_M2 5000_2000_M2 0.015
r 5000_2000_M2 5000_3000_M2 0.015
r 5000_3000_M2 5000_4000_M2 0.015
r 5000_4000_M2 5000_5000_M2 0.015

* ============================================================================
* Via connections (M1 to M2) at each grid point
* ============================================================================

* Via resistance: 0.005 Ohm per via
r 1000_1000_M1 1000_1000_M2 0.005
r 2000_1000_M1 2000_1000_M2 0.005
r 3000_1000_M1 3000_1000_M2 0.005
r 4000_1000_M1 4000_1000_M2 0.005
r 5000_1000_M1 5000_1000_M2 0.005

r 1000_2000_M1 1000_2000_M2 0.005
r 2000_2000_M1 2000_2000_M2 0.005
r 3000_2000_M1 3000_2000_M2 0.005
r 4000_2000_M1 4000_2000_M2 0.005
r 5000_2000_M1 5000_2000_M2 0.005

r 1000_3000_M1 1000_3000_M2 0.005
r 2000_3000_M1 2000_3000_M2 0.005
r 3000_3000_M1 3000_3000_M2 0.005
r 4000_3000_M1 4000_3000_M2 0.005
r 5000_3000_M1 5000_3000_M2 0.005

r 1000_4000_M1 1000_4000_M2 0.005
r 2000_4000_M1 2000_4000_M2 0.005
r 3000_4000_M1 3000_4000_M2 0.005
r 4000_4000_M1 4000_4000_M2 0.005
r 5000_4000_M1 5000_4000_M2 0.005

r 1000_5000_M1 1000_5000_M2 0.005
r 2000_5000_M1 2000_5000_M2 0.005
r 3000_5000_M1 3000_5000_M2 0.005
r 4000_5000_M1 4000_5000_M2 0.005
r 5000_5000_M1 5000_5000_M2 0.005

* ============================================================================
* Decoupling capacitors to ground (every grid point on both layers)
* ============================================================================

* M1 layer capacitors (1 pF each)
c 1000_1000_M1 0 1e-12
c 2000_1000_M1 0 1e-12
c 3000_1000_M1 0 1e-12
c 4000_1000_M1 0 1e-12
c 5000_1000_M1 0 1e-12

c 1000_2000_M1 0 1e-12
c 2000_2000_M1 0 1e-12
c 3000_2000_M1 0 1e-12
c 4000_2000_M1 0 1e-12
c 5000_2000_M1 0 1e-12

c 1000_3000_M1 0 1e-12
c 2000_3000_M1 0 1e-12
c 3000_3000_M1 0 1e-12
c 4000_3000_M1 0 1e-12
c 5000_3000_M1 0 1e-12

c 1000_4000_M1 0 1e-12
c 2000_4000_M1 0 1e-12
c 3000_4000_M1 0 1e-12
c 4000_4000_M1 0 1e-12
c 5000_4000_M1 0 1e-12

c 1000_5000_M1 0 1e-12
c 2000_5000_M1 0 1e-12
c 3000_5000_M1 0 1e-12
c 4000_5000_M1 0 1e-12
c 5000_5000_M1 0 1e-12

* M2 layer capacitors (1 pF each)
c 1000_1000_M2 0 1e-12
c 2000_1000_M2 0 1e-12
c 3000_1000_M2 0 1e-12
c 4000_1000_M2 0 1e-12
c 5000_1000_M2 0 1e-12

c 1000_2000_M2 0 1e-12
c 2000_2000_M2 0 1e-12
c 3000_2000_M2 0 1e-12
c 4000_2000_M2 0 1e-12
c 5000_2000_M2 0 1e-12

c 1000_3000_M2 0 1e-12
c 2000_3000_M2 0 1e-12
c 3000_3000_M2 0 1e-12
c 4000_3000_M2 0 1e-12
c 5000_3000_M2 0 1e-12

c 1000_4000_M2 0 1e-12
c 2000_4000_M2 0 1e-12
c 3000_4000_M2 0 1e-12
c 4000_4000_M2 0 1e-12
c 5000_4000_M2 0 1e-12

c 1000_5000_M2 0 1e-12
c 2000_5000_M2 0 1e-12
c 3000_5000_M2 0 1e-12
c 4000_5000_M2 0 1e-12
c 5000_5000_M2 0 1e-12
